//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT103), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G8gat), .B(G36gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(KEYINPUT86), .B(new_n213_), .C1(new_n214_), .C2(new_n212_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT22), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G169gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n217_), .A2(new_n212_), .A3(KEYINPUT86), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(G176gat), .B1(new_n215_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n209_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT23), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n216_), .A2(G169gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n210_), .A2(KEYINPUT22), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT85), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n218_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT87), .B(new_n223_), .C1(new_n234_), .C2(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n225_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G197gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT21), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G211gat), .B(G218gat), .Z(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(KEYINPUT21), .C1(new_n241_), .C2(new_n243_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n210_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT24), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n254_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT26), .B(G190gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT25), .B1(new_n254_), .B2(KEYINPUT82), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n253_), .A2(KEYINPUT84), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT84), .B1(new_n253_), .B2(new_n258_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n227_), .B(new_n252_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n236_), .A2(new_n249_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT100), .B1(new_n229_), .B2(new_n230_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT100), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n211_), .A2(new_n217_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(G176gat), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT101), .B1(new_n266_), .B2(new_n224_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n211_), .A2(new_n217_), .A3(new_n264_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n250_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT101), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n223_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n228_), .A3(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(new_n251_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT25), .B(G183gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n256_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n221_), .A3(new_n251_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n275_), .A2(new_n227_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n249_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n262_), .A2(new_n282_), .A3(KEYINPUT20), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n236_), .A2(new_n261_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n281_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n285_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n273_), .A2(new_n249_), .A3(new_n279_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n288_), .A2(KEYINPUT20), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT102), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT102), .B1(new_n283_), .B2(new_n285_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n208_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT102), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n298_), .A2(new_n207_), .A3(new_n294_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n202_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(new_n208_), .A3(new_n295_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n288_), .A2(KEYINPUT20), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n289_), .B1(new_n302_), .B2(new_n290_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n283_), .A2(new_n285_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n207_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(KEYINPUT27), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT92), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n314_));
  OR2_X1    g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT92), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n323_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n335_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n314_), .A2(new_n316_), .A3(new_n315_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n316_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n312_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n322_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n331_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n334_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n323_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n346_), .A2(KEYINPUT104), .A3(KEYINPUT4), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n335_), .A2(new_n336_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n349_), .A3(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT104), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n348_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n339_), .B1(new_n354_), .B2(new_n338_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  INV_X1    g155(.A(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n355_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n300_), .A2(new_n306_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT28), .B(G22gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n344_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n368_));
  INV_X1    g167(.A(G50gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n330_), .A2(new_n315_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n311_), .A2(new_n370_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(G50gat), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n369_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n366_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT94), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT97), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT93), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n281_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n372_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  NOR4_X1   g186(.A1(new_n386_), .A2(KEYINPUT93), .A3(new_n387_), .A4(new_n249_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n382_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT93), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n281_), .B(new_n390_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n393_), .A2(new_n390_), .A3(new_n383_), .A4(new_n281_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n394_), .C1(KEYINPUT97), .C2(new_n381_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n379_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n381_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n392_), .A2(KEYINPUT95), .A3(new_n397_), .A4(new_n394_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n398_), .A2(new_n378_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n381_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n399_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n400_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n396_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT98), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n402_), .A2(new_n381_), .A3(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(new_n378_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT96), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n399_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n396_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n236_), .A2(new_n416_), .A3(new_n261_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n236_), .B2(new_n261_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT90), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n287_), .A2(KEYINPUT30), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n417_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G71gat), .B(G99gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT89), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT88), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n427_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n420_), .A2(new_n423_), .A3(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n421_), .A2(new_n430_), .A3(new_n422_), .A4(new_n417_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT91), .A3(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n334_), .B(KEYINPUT31), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(KEYINPUT91), .A3(new_n433_), .A4(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n408_), .A2(new_n415_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n365_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n414_), .B1(new_n413_), .B2(new_n396_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n396_), .ZN(new_n444_));
  AOI211_X1 g243(.A(KEYINPUT98), .B(new_n444_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT33), .B1(new_n355_), .B2(new_n361_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n346_), .A2(KEYINPUT4), .A3(new_n347_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT104), .B1(new_n336_), .B2(new_n349_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n337_), .B1(new_n450_), .B2(new_n348_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  NOR4_X1   g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n339_), .A4(new_n360_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n207_), .B1(new_n298_), .B2(new_n294_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n338_), .B1(new_n450_), .B2(new_n348_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT105), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n346_), .A2(new_n338_), .A3(new_n347_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(KEYINPUT105), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n457_), .A2(new_n360_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n301_), .A2(new_n454_), .A3(new_n455_), .A4(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n208_), .A2(KEYINPUT32), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n293_), .A2(new_n295_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n362_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n439_), .B1(new_n461_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n446_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n442_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G230gat), .ZN(new_n470_));
  INV_X1    g269(.A(G233gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT65), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G85gat), .B(G92gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT9), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n357_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n357_), .A2(KEYINPUT64), .ZN(new_n487_));
  OAI21_X1  g286(.A(G92gat), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT10), .B(G99gat), .Z(new_n489_));
  INV_X1    g288(.A(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n482_), .A2(new_n485_), .A3(new_n488_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n494_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT67), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n496_), .B2(KEYINPUT7), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  OAI221_X1 g297(.A(new_n494_), .B1(G99gat), .B2(G106gat), .C1(new_n496_), .C2(KEYINPUT7), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n478_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT69), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT69), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(new_n503_), .A3(new_n484_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(KEYINPUT8), .A3(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n498_), .A2(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n482_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n484_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n493_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n473_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n500_), .A2(new_n503_), .A3(new_n484_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n503_), .B1(new_n500_), .B2(new_n484_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  AOI211_X1 g322(.A(new_n483_), .B(new_n508_), .C1(new_n482_), .C2(new_n506_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n492_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n473_), .A3(new_n526_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n472_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(KEYINPUT70), .A3(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n511_), .A2(new_n518_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n472_), .B(new_n532_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G176gat), .B(G204gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n531_), .A2(new_n536_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n536_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(new_n530_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT72), .B(new_n541_), .C1(new_n544_), .C2(new_n530_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT73), .B(G29gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(G43gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n369_), .ZN(new_n561_));
  INV_X1    g360(.A(G36gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n559_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G36gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n558_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G1gat), .B(G8gat), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n575_));
  INV_X1    g374(.A(G1gat), .ZN(new_n576_));
  INV_X1    g375(.A(G8gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n575_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n573_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT77), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n572_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n571_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n571_), .A2(new_n581_), .A3(new_n585_), .A4(KEYINPUT78), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n571_), .B1(new_n585_), .B2(new_n581_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT79), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT79), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n594_), .B(new_n591_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n557_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n571_), .B(KEYINPUT15), .ZN(new_n597_));
  INV_X1    g396(.A(new_n585_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n581_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n556_), .A3(new_n590_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n555_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n601_), .A3(new_n555_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT80), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT81), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT81), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n602_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n469_), .A2(new_n551_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT76), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(KEYINPUT76), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT34), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n525_), .A2(new_n597_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT74), .ZN(new_n629_));
  INV_X1    g428(.A(new_n571_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n525_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n511_), .A2(KEYINPUT74), .A3(new_n571_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n627_), .A2(new_n624_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n628_), .A2(new_n631_), .A3(new_n636_), .A4(new_n632_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n623_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT75), .B1(new_n635_), .B2(new_n637_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  AOI221_X4 g441(.A(KEYINPUT75), .B1(new_n642_), .B2(new_n623_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n617_), .B(new_n618_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(new_n640_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n643_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(KEYINPUT76), .A3(new_n616_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n644_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n518_), .B(new_n651_), .Z(new_n652_));
  NOR2_X1   g451(.A1(new_n599_), .A2(new_n598_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT17), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(G211gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G183gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  NOR3_X1   g458(.A1(new_n654_), .A2(new_n655_), .A3(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(KEYINPUT17), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n654_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n650_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n615_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n576_), .A3(new_n362_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT38), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n641_), .A2(new_n643_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n663_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n615_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n363_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n673_), .ZN(G1324gat));
  NAND2_X1  g473(.A1(new_n300_), .A2(new_n306_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G8gat), .B1(new_n672_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT39), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n666_), .A2(new_n577_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  INV_X1    g481(.A(new_n439_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G15gat), .B1(new_n672_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT41), .Z(new_n685_));
  NOR3_X1   g484(.A1(new_n665_), .A2(G15gat), .A3(new_n683_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT106), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1326gat));
  OAI21_X1  g487(.A(G22gat), .B1(new_n672_), .B2(new_n446_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT42), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n446_), .A2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n665_), .B2(new_n691_), .ZN(G1327gat));
  NAND3_X1  g491(.A1(new_n551_), .A2(new_n663_), .A3(new_n614_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n669_), .B1(new_n442_), .B2(new_n468_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n362_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n469_), .B2(new_n650_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n683_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n408_), .A2(new_n415_), .A3(new_n439_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n364_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n446_), .A2(new_n467_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n698_), .B(new_n650_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n694_), .B1(new_n699_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(KEYINPUT107), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n650_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT43), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n693_), .B1(new_n711_), .B2(new_n704_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(G29gat), .A3(new_n362_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT44), .B(new_n694_), .C1(new_n699_), .C2(new_n705_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT108), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n697_), .B1(new_n715_), .B2(new_n721_), .ZN(G1328gat));
  OAI21_X1  g521(.A(new_n675_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n706_), .B2(new_n707_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n712_), .A2(new_n709_), .A3(KEYINPUT44), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G36gat), .B1(new_n723_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n696_), .A2(new_n562_), .A3(new_n675_), .ZN(new_n730_));
  XOR2_X1   g529(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .A4(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n728_), .A2(new_n729_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n716_), .A2(new_n717_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n712_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n676_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n562_), .B1(new_n738_), .B2(new_n714_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n732_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n734_), .B(new_n735_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n733_), .A2(new_n741_), .ZN(G1329gat));
  INV_X1    g541(.A(new_n696_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n560_), .B1(new_n743_), .B2(new_n683_), .ZN(new_n744_));
  OAI211_X1 g543(.A(G43gat), .B(new_n439_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n726_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g546(.A(new_n369_), .B1(new_n743_), .B2(new_n446_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n446_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n714_), .A2(G50gat), .A3(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(new_n720_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT111), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n748_), .C1(new_n750_), .C2(new_n720_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1331gat));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n614_), .B(new_n551_), .C1(new_n442_), .C2(new_n468_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n664_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n758_), .B2(new_n363_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT112), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n671_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n362_), .A2(G57gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT113), .ZN(G1332gat));
  OAI21_X1  g563(.A(G64gat), .B1(new_n761_), .B2(new_n676_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT48), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n676_), .A2(G64gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n758_), .B2(new_n767_), .ZN(G1333gat));
  OAI21_X1  g567(.A(G71gat), .B1(new_n761_), .B2(new_n683_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT49), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n683_), .A2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n758_), .B2(new_n771_), .ZN(G1334gat));
  OAI21_X1  g571(.A(G78gat), .B1(new_n761_), .B2(new_n446_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT50), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n446_), .A2(G78gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n758_), .B2(new_n775_), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n551_), .A2(new_n662_), .A3(new_n614_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n695_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n362_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n777_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n711_), .B2(new_n704_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n357_), .A2(KEYINPUT64), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n362_), .B1(new_n487_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT114), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(new_n782_), .B2(new_n785_), .ZN(G1336gat));
  AOI21_X1  g585(.A(G92gat), .B1(new_n779_), .B2(new_n675_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n675_), .A2(G92gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n782_), .B2(new_n788_), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n489_), .A3(new_n439_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT115), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n782_), .A2(new_n439_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(G99gat), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n779_), .A2(new_n490_), .A3(new_n749_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n490_), .B1(new_n782_), .B2(new_n749_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n798_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g601(.A1(new_n644_), .A2(new_n649_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n528_), .A2(new_n529_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n472_), .ZN(new_n805_));
  AND2_X1   g604(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n528_), .A2(new_n472_), .A3(new_n529_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n806_), .B1(new_n530_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n541_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT56), .B(new_n541_), .C1(new_n809_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n556_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n600_), .A2(new_n557_), .A3(new_n590_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n554_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n604_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n543_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n543_), .A3(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT58), .B1(new_n817_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n803_), .B2(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n815_), .A2(new_n816_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT58), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n650_), .B(new_n831_), .C1(new_n829_), .C2(KEYINPUT58), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n543_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n817_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n547_), .A2(new_n548_), .A3(new_n821_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  INV_X1    g640(.A(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n817_), .B2(new_n836_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n670_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n663_), .B1(new_n834_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n614_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n664_), .A2(new_n551_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n850_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n664_), .A2(new_n551_), .A3(new_n847_), .A4(new_n851_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n846_), .A2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(new_n362_), .A3(new_n440_), .A4(new_n676_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n614_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n675_), .B1(new_n846_), .B2(new_n856_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT59), .A3(new_n362_), .A4(new_n440_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n669_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n843_), .A2(new_n841_), .A3(new_n670_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n662_), .B1(new_n866_), .B2(new_n833_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n855_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n362_), .B(new_n676_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n869_), .B2(new_n701_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n847_), .B1(new_n862_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n860_), .B1(new_n871_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n551_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n859_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n873_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n551_), .B1(new_n862_), .B2(new_n870_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n873_), .ZN(G1341gat));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n858_), .B2(new_n663_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT120), .B(new_n878_), .C1(new_n858_), .C2(new_n663_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n862_), .A2(new_n870_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n662_), .A2(G127gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT121), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n881_), .A2(new_n882_), .B1(new_n883_), .B2(new_n885_), .ZN(G1342gat));
  NOR3_X1   g685(.A1(new_n869_), .A2(new_n669_), .A3(new_n701_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n887_), .B2(G134gat), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n889_), .B(new_n890_), .C1(new_n858_), .C2(new_n669_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT123), .B(G134gat), .Z(new_n893_));
  AOI211_X1 g692(.A(new_n803_), .B(new_n893_), .C1(new_n862_), .C2(new_n870_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n869_), .A2(new_n700_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n614_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g697(.A(new_n551_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n662_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  AOI21_X1  g703(.A(G162gat), .B1(new_n896_), .B2(new_n670_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n650_), .A2(G162gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n896_), .B2(new_n906_), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n676_), .A2(new_n362_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n440_), .B(new_n908_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909_), .B2(new_n847_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n913_), .B(G169gat), .C1(new_n909_), .C2(new_n847_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n912_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(KEYINPUT125), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n268_), .A2(new_n269_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n909_), .A2(new_n847_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(new_n917_), .C1(new_n918_), .C2(new_n919_), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n909_), .A2(new_n551_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n250_), .ZN(G1349gat));
  NOR2_X1   g721(.A1(new_n909_), .A2(new_n663_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n276_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n254_), .B2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n909_), .B2(new_n803_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n670_), .A2(new_n256_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n909_), .B2(new_n927_), .ZN(G1351gat));
  AND2_X1   g727(.A1(new_n857_), .A2(new_n908_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n441_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n240_), .A3(new_n614_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G197gat), .B1(new_n930_), .B2(new_n847_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n242_), .A2(KEYINPUT126), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n242_), .A2(KEYINPUT126), .ZN(new_n936_));
  OAI22_X1  g735(.A1(new_n930_), .A2(new_n551_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n931_), .A2(new_n899_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n935_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n930_), .B2(new_n663_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  NAND4_X1  g741(.A1(new_n929_), .A2(new_n662_), .A3(new_n441_), .A4(new_n942_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1354gat));
  NAND2_X1  g743(.A1(new_n650_), .A2(G218gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT127), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n929_), .A2(new_n670_), .A3(new_n441_), .ZN(new_n947_));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  AOI22_X1  g747(.A1(new_n931_), .A2(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1355gat));
endmodule


