//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  NOR2_X1   g000(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n212_), .B(G85gat), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n215_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(G106gat), .B1(new_n206_), .B2(new_n208_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NOR3_X1   g032(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n231_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n210_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(KEYINPUT68), .A3(new_n232_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n223_), .A3(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n216_), .A2(new_n217_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n230_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n230_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n220_), .A2(new_n222_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n232_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n223_), .A2(new_n247_), .A3(new_n238_), .A4(new_n232_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  OAI22_X1  g048(.A1(new_n225_), .A2(new_n229_), .B1(new_n242_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G29gat), .B(G36gat), .Z(new_n251_));
  XOR2_X1   g050(.A(G43gat), .B(G50gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G29gat), .B(G36gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT35), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n250_), .A2(new_n259_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265_));
  INV_X1    g064(.A(new_n257_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n250_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n240_), .A2(new_n241_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT8), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n246_), .A2(new_n248_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n243_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n228_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n211_), .A2(KEYINPUT66), .A3(new_n224_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n269_), .A2(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT74), .A3(new_n257_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n267_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n263_), .A2(new_n260_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n264_), .A2(new_n267_), .A3(new_n276_), .A4(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G190gat), .B(G218gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT75), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT36), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n285_), .B(KEYINPUT36), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT37), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT76), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(KEYINPUT37), .C1(new_n288_), .C2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n279_), .A2(new_n281_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n289_), .B1(new_n295_), .B2(KEYINPUT77), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n279_), .A2(new_n297_), .A3(new_n281_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n288_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT37), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n292_), .A2(new_n294_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(KEYINPUT78), .A2(G15gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT78), .A2(G15gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(G22gat), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(G22gat), .B1(new_n305_), .B2(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n304_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n309_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n307_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n304_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G64gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n319_));
  XOR2_X1   g118(.A(G71gat), .B(G78gat), .Z(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G231gat), .ZN(new_n328_));
  INV_X1    g127(.A(G233gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n317_), .A2(new_n325_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G127gat), .B(G155gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G183gat), .B(G211gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT17), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n332_), .A2(new_n343_), .A3(new_n333_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n301_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G120gat), .B(G148gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n353_), .A2(KEYINPUT72), .A3(new_n354_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G230gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n325_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n275_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n275_), .A2(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n361_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n275_), .B2(new_n362_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n361_), .B1(new_n275_), .B2(new_n362_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n250_), .A2(KEYINPUT12), .A3(new_n325_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n359_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n366_), .A2(new_n371_), .A3(new_n355_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT13), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT13), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G113gat), .B(G141gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G169gat), .B(G197gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n315_), .B1(new_n314_), .B2(new_n304_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n304_), .ZN(new_n385_));
  AOI211_X1 g184(.A(new_n311_), .B(new_n385_), .C1(new_n313_), .C2(new_n307_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n253_), .A2(KEYINPUT80), .A3(new_n256_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT80), .B1(new_n253_), .B2(new_n256_), .ZN(new_n389_));
  OAI22_X1  g188(.A1(new_n384_), .A2(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n257_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n312_), .A2(new_n392_), .A3(new_n316_), .A4(new_n387_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT81), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT81), .B1(new_n390_), .B2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G229gat), .A2(G233gat), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n259_), .A2(new_n317_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n396_), .A3(new_n393_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n383_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n395_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n396_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT81), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n399_), .A3(new_n382_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n379_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(G190gat), .ZN(new_n414_));
  INV_X1    g213(.A(G190gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT25), .B(G183gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT83), .B(KEYINPUT26), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(new_n415_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT23), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(G183gat), .A3(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n432_));
  INV_X1    g231(.A(G183gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n415_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n421_), .A2(new_n423_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT85), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n441_), .A2(new_n442_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n440_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n439_), .A3(new_n443_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n431_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT30), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT86), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G43gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(G15gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n452_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n449_), .A2(KEYINPUT86), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n456_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461_));
  INV_X1    g260(.A(G120gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G113gat), .ZN(new_n463_));
  INV_X1    g262(.A(G113gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G120gat), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT87), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT87), .B1(new_n463_), .B2(new_n465_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n461_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n464_), .A2(G120gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n462_), .A2(G113gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT87), .ZN(new_n473_));
  XOR2_X1   g272(.A(G127gat), .B(G134gat), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT88), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n458_), .A2(new_n460_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n449_), .A2(KEYINPUT86), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n456_), .B1(new_n485_), .B2(new_n459_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n460_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G228gat), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n490_), .A2(new_n329_), .A3(KEYINPUT92), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G197gat), .A2(G204gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT21), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT21), .ZN(new_n497_));
  AND2_X1   g296(.A1(G197gat), .A2(G204gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n493_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G211gat), .B(G218gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G218gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G211gat), .ZN(new_n503_));
  INV_X1    g302(.A(G211gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G218gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(KEYINPUT21), .A3(new_n494_), .A4(new_n495_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G141gat), .ZN(new_n509_));
  INV_X1    g308(.A(G148gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(KEYINPUT3), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT3), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(G141gat), .B2(G148gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G141gat), .A2(G148gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT2), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT90), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n514_), .A2(new_n517_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G155gat), .B(G162gat), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT1), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n509_), .A2(new_n510_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n526_), .A2(new_n515_), .A3(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n522_), .A2(new_n523_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n508_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT92), .B1(new_n490_), .B2(new_n329_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G78gat), .B(G106gat), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n492_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n522_), .A2(new_n523_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n525_), .A2(new_n528_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n530_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n501_), .A2(new_n507_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n532_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n491_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n545_), .A3(KEYINPUT91), .ZN(new_n546_));
  INV_X1    g345(.A(new_n529_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT28), .B1(new_n547_), .B2(KEYINPUT29), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n529_), .A2(new_n549_), .A3(new_n530_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G22gat), .B(G50gat), .Z(new_n551_));
  AND3_X1   g350(.A1(new_n548_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n553_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n556_), .A2(new_n536_), .A3(new_n545_), .A4(KEYINPUT91), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n480_), .A2(new_n547_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G225gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n466_), .A2(new_n467_), .A3(new_n461_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n478_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n468_), .A2(new_n475_), .A3(KEYINPUT95), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n529_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G29gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G85gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT0), .B(G57gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT4), .B1(new_n480_), .B2(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n559_), .A2(new_n565_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n573_), .B2(KEYINPUT4), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n560_), .B(KEYINPUT96), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n566_), .B(new_n571_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT4), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n575_), .B1(new_n581_), .B2(new_n572_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(KEYINPUT33), .A3(new_n566_), .A4(new_n571_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G226gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT19), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT93), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n540_), .A2(new_n431_), .A3(new_n447_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT26), .B(G190gat), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n418_), .A2(new_n588_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n429_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT22), .B(G169gat), .ZN(new_n591_));
  INV_X1    g390(.A(G176gat), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n425_), .A2(new_n434_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n589_), .A2(new_n430_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT20), .B1(new_n595_), .B2(new_n540_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n586_), .B1(new_n587_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n448_), .A2(new_n508_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n585_), .B1(new_n595_), .B2(new_n540_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT20), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G8gat), .B(G36gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G64gat), .B(G92gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n605_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n597_), .A2(new_n610_), .A3(new_n600_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n560_), .ZN(new_n613_));
  OAI221_X1 g412(.A(new_n570_), .B1(new_n573_), .B2(new_n576_), .C1(new_n574_), .C2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n579_), .A2(new_n583_), .A3(new_n612_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n597_), .A2(new_n600_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT20), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n593_), .A2(new_n594_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n415_), .A2(KEYINPUT26), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n433_), .A2(KEYINPUT25), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G183gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n413_), .A2(G190gat), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .A4(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n430_), .A2(new_n425_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n618_), .B1(new_n627_), .B2(new_n508_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n540_), .A2(new_n431_), .A3(new_n447_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n586_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n598_), .A2(KEYINPUT20), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n619_), .A2(new_n626_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n508_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n585_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n617_), .A2(new_n632_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n610_), .A2(KEYINPUT32), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n618_), .B1(new_n448_), .B2(new_n508_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n586_), .A2(new_n630_), .B1(new_n643_), .B2(new_n599_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n640_), .A3(KEYINPUT97), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n582_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n571_), .B1(new_n582_), .B2(new_n566_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n642_), .B(new_n645_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n558_), .B1(new_n615_), .B2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n609_), .A2(new_n611_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT27), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n644_), .B2(new_n610_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n585_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n636_), .A2(new_n508_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n635_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n654_), .B1(new_n657_), .B2(new_n643_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n608_), .B1(new_n658_), .B2(new_n631_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n651_), .A2(new_n652_), .B1(new_n653_), .B2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n650_), .A2(new_n558_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n489_), .B1(new_n649_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n660_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n558_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n483_), .A2(new_n488_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n650_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n411_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n346_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n650_), .B(KEYINPUT99), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n302_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT38), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n299_), .B(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n662_), .A2(new_n666_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n650_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n411_), .A2(new_n345_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n671_), .B1(new_n681_), .B2(new_n302_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT102), .Z(G1324gat));
  NAND3_X1  g482(.A1(new_n668_), .A2(new_n303_), .A3(new_n663_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n677_), .A2(new_n663_), .A3(new_n679_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G8gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G8gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  NAND3_X1  g490(.A1(new_n668_), .A2(new_n454_), .A3(new_n665_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n677_), .A2(new_n665_), .A3(new_n679_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(new_n693_), .B2(G15gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n668_), .A2(new_n697_), .A3(new_n558_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n677_), .A2(new_n558_), .A3(new_n679_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(G22gat), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(new_n299_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n345_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n667_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n678_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n411_), .A2(new_n705_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n674_), .A2(new_n711_), .A3(new_n301_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n674_), .B2(new_n301_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n710_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716_));
  INV_X1    g515(.A(new_n710_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n674_), .A2(new_n301_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT43), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n674_), .A2(new_n301_), .A3(new_n711_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n721_), .B2(KEYINPUT44), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(KEYINPUT104), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n715_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(KEYINPUT105), .A3(new_n669_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n726_), .B2(new_n669_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n709_), .B1(new_n728_), .B2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n733_));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n726_), .B2(new_n663_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n707_), .A2(new_n734_), .A3(new_n663_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n736_), .B(new_n737_), .Z(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n732_), .B(new_n733_), .C1(new_n735_), .C2(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n721_), .A2(new_n716_), .A3(KEYINPUT44), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT104), .B1(new_n723_), .B2(new_n724_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n663_), .B(new_n714_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G36gat), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n744_), .A2(KEYINPUT107), .A3(new_n731_), .A4(new_n738_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n740_), .A2(new_n745_), .ZN(G1329gat));
  AOI21_X1  g545(.A(G43gat), .B1(new_n707_), .B2(new_n665_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n665_), .A2(G43gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n726_), .B2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g549(.A(G50gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n707_), .A2(new_n751_), .A3(new_n558_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n714_), .A2(new_n558_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n753_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT108), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n756_), .A2(KEYINPUT109), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT109), .B1(new_n756_), .B2(new_n759_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n752_), .B1(new_n760_), .B2(new_n761_), .ZN(G1331gat));
  NOR3_X1   g561(.A1(new_n379_), .A2(new_n410_), .A3(new_n345_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n677_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n677_), .A2(KEYINPUT110), .A3(new_n763_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(G57gat), .A3(new_n678_), .A4(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n379_), .A2(new_n410_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n674_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n346_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G57gat), .B1(new_n774_), .B2(new_n669_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n769_), .A2(new_n770_), .A3(new_n775_), .ZN(G1332gat));
  OR3_X1    g575(.A1(new_n773_), .A2(G64gat), .A3(new_n660_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n663_), .A3(new_n767_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(G64gat), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G64gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1333gat));
  OR3_X1    g581(.A1(new_n773_), .A2(G71gat), .A3(new_n489_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n766_), .A2(new_n665_), .A3(new_n767_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(G71gat), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G71gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  INV_X1    g587(.A(new_n558_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n773_), .A2(G78gat), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n766_), .A2(new_n558_), .A3(new_n767_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(G78gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n791_), .B2(G78gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1335gat));
  AND2_X1   g594(.A1(new_n772_), .A2(new_n706_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n669_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n771_), .A2(new_n345_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n678_), .A2(G85gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT114), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n797_), .B1(new_n799_), .B2(new_n801_), .ZN(G1336gat));
  AOI21_X1  g601(.A(G92gat), .B1(new_n796_), .B2(new_n663_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n213_), .A2(new_n214_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n660_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n803_), .B1(new_n799_), .B2(new_n805_), .ZN(G1337gat));
  AOI21_X1  g605(.A(new_n237_), .B1(new_n799_), .B2(new_n665_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n665_), .A2(new_n209_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n796_), .B2(new_n808_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g609(.A1(new_n796_), .A2(new_n210_), .A3(new_n558_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n799_), .A2(new_n558_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n210_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g617(.A1(new_n345_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n373_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n377_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n379_), .A2(KEYINPUT116), .A3(new_n819_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n292_), .A2(new_n294_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT37), .B2(new_n704_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n357_), .A2(new_n358_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n368_), .A2(new_n363_), .A3(new_n370_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n834_), .A2(new_n371_), .B1(new_n835_), .B2(new_n361_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n368_), .A2(new_n369_), .A3(KEYINPUT55), .A4(new_n370_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n371_), .A2(new_n834_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n361_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n837_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n359_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT56), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n403_), .A2(new_n396_), .A3(new_n405_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n393_), .A2(new_n404_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n382_), .B1(new_n847_), .B2(new_n398_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n374_), .A2(new_n407_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n840_), .A2(new_n845_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n840_), .A2(new_n845_), .A3(KEYINPUT58), .A4(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n301_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n375_), .A2(new_n407_), .A3(new_n849_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n366_), .A2(new_n371_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n857_), .A2(new_n355_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n838_), .B2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n844_), .A2(new_n859_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n704_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(new_n704_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n855_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n705_), .B1(new_n867_), .B2(KEYINPUT118), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n855_), .B(new_n869_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n832_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n669_), .A2(new_n665_), .A3(new_n664_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n464_), .A3(new_n410_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n867_), .A2(new_n345_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n875_), .A2(new_n832_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  INV_X1    g676(.A(new_n872_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(new_n410_), .C1(new_n877_), .C2(new_n873_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n874_), .B1(new_n881_), .B2(new_n464_), .ZN(G1340gat));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G120gat), .B1(new_n883_), .B2(new_n379_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n873_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n462_), .B1(new_n379_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(KEYINPUT60), .B2(new_n462_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n885_), .B2(new_n887_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n873_), .A2(new_n889_), .A3(new_n705_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n879_), .B(new_n705_), .C1(new_n877_), .C2(new_n873_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n892_), .B2(new_n889_), .ZN(G1342gat));
  NAND2_X1  g692(.A1(new_n301_), .A2(G134gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT119), .Z(new_n895_));
  OAI211_X1 g694(.A(new_n879_), .B(new_n895_), .C1(new_n877_), .C2(new_n873_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n673_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G134gat), .B1(new_n873_), .B2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1343gat));
  NAND4_X1  g699(.A1(new_n669_), .A2(new_n489_), .A3(new_n558_), .A4(new_n660_), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT120), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n871_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n410_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g704(.A(new_n379_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n705_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  NOR4_X1   g710(.A1(new_n871_), .A2(G162gat), .A3(new_n673_), .A4(new_n902_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914_));
  INV_X1    g713(.A(G162gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n871_), .A2(new_n828_), .A3(new_n902_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n913_), .B(new_n914_), .C1(new_n915_), .C2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n915_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n918_), .B2(new_n912_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1347gat));
  INV_X1    g719(.A(new_n669_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n665_), .A3(new_n663_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n789_), .B(new_n923_), .C1(new_n875_), .C2(new_n832_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924_), .B2(new_n409_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n926_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n924_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n929_), .A2(new_n591_), .A3(new_n410_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(G1348gat));
  OAI21_X1  g730(.A(new_n592_), .B1(new_n924_), .B2(new_n379_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n867_), .A2(KEYINPUT118), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n934_), .A2(new_n345_), .A3(new_n870_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n832_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n558_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n923_), .A2(G176gat), .A3(new_n906_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n933_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n558_), .A4(new_n938_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n932_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT123), .B(new_n932_), .C1(new_n940_), .C2(new_n941_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n876_), .A2(new_n789_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n923_), .A2(new_n705_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n947_), .A2(new_n418_), .A3(new_n948_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n871_), .A2(new_n558_), .A3(new_n948_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n950_), .A2(KEYINPUT124), .ZN(new_n951_));
  AOI21_X1  g750(.A(G183gat), .B1(new_n950_), .B2(KEYINPUT124), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n951_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n924_), .B2(new_n828_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n898_), .A2(new_n588_), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n955_), .B(KEYINPUT125), .Z(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n924_), .B2(new_n956_), .ZN(G1351gat));
  NAND2_X1  g756(.A1(new_n935_), .A2(new_n936_), .ZN(new_n958_));
  NOR4_X1   g757(.A1(new_n665_), .A2(new_n678_), .A3(new_n789_), .A4(new_n660_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n409_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT126), .B(G197gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1352gat));
  INV_X1    g762(.A(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n906_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g765(.A(new_n345_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n964_), .A2(new_n968_), .ZN(new_n969_));
  OR2_X1    g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n960_), .B2(new_n828_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n898_), .A2(new_n502_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n960_), .B2(new_n973_), .ZN(G1355gat));
endmodule


