//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT12), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n213_), .B(new_n214_), .C1(new_n215_), .C2(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  XOR2_X1   g025(.A(G85gat), .B(G92gat), .Z(new_n227_));
  AND3_X1   g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n219_), .A2(KEYINPUT66), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n216_), .A2(new_n218_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n224_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n227_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n230_), .B1(new_n235_), .B2(KEYINPUT8), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT67), .B(new_n226_), .C1(new_n234_), .C2(new_n227_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT68), .ZN(new_n239_));
  INV_X1    g038(.A(new_n227_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n219_), .A2(KEYINPUT66), .B1(new_n221_), .B2(new_n223_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n233_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n226_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n216_), .A2(new_n218_), .A3(new_n232_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n232_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n224_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n230_), .B(KEYINPUT8), .C1(new_n247_), .C2(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n229_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n239_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n240_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT10), .B(G99gat), .Z(new_n257_));
  AOI21_X1  g056(.A(new_n246_), .B1(new_n214_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n212_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n250_), .B1(new_n249_), .B2(new_n229_), .ZN(new_n261_));
  AOI211_X1 g060(.A(KEYINPUT68), .B(new_n228_), .C1(new_n243_), .C2(new_n248_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n212_), .B(new_n259_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n211_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n238_), .A2(new_n208_), .A3(new_n259_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G230gat), .A2(G233gat), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n266_), .A2(KEYINPUT70), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT70), .B1(new_n266_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n238_), .A2(new_n259_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n209_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT12), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n267_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n266_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G120gat), .B(G148gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G176gat), .B(G204gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT72), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT72), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n277_), .A2(new_n280_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n285_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(KEYINPUT13), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT13), .B1(new_n290_), .B2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT103), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT85), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n300_), .B(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT81), .B(G190gat), .Z(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(KEYINPUT26), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT25), .B(G183gat), .Z(new_n314_));
  OAI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G183gat), .A3(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT23), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n317_), .A2(new_n318_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n316_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n320_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n312_), .B2(G183gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G169gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G15gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  INV_X1    g138(.A(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n338_), .B(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n305_), .B1(new_n344_), .B2(KEYINPUT87), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(KEYINPUT87), .B2(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(KEYINPUT87), .A3(new_n305_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT90), .B(G197gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  INV_X1    g150(.A(G204gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT92), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G211gat), .B(G218gat), .Z(new_n359_));
  OR2_X1    g158(.A1(new_n349_), .A2(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(G197gat), .B2(G204gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n353_), .A4(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G141gat), .ZN(new_n372_));
  INV_X1    g171(.A(G148gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT3), .ZN(new_n375_));
  OR3_X1    g174(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(new_n376_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT88), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n369_), .B(new_n371_), .C1(new_n379_), .C2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n370_), .B1(KEYINPUT1), .B2(new_n369_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(KEYINPUT1), .B2(new_n369_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n378_), .A3(new_n374_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n366_), .B(new_n367_), .C1(new_n368_), .C2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n368_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT93), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n366_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n364_), .A2(KEYINPUT93), .A3(new_n365_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n392_), .B2(new_n367_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G78gat), .B(G106gat), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n386_), .A2(new_n368_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n394_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n387_), .C1(new_n392_), .C2(new_n367_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n395_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G57gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n386_), .B1(new_n302_), .B2(new_n299_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n386_), .B2(new_n303_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT100), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(KEYINPUT100), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n303_), .A2(new_n386_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT4), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n412_), .B2(KEYINPUT4), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n415_), .B(new_n416_), .C1(new_n417_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(new_n413_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n409_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT26), .B(G190gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT94), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n310_), .B1(new_n432_), .B2(new_n314_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n318_), .B1(new_n325_), .B2(new_n320_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n333_), .B1(new_n326_), .B2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n439_), .B(KEYINPUT96), .Z(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n430_), .B1(new_n441_), .B2(new_n366_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n366_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(new_n334_), .A3(new_n329_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT19), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT18), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G64gat), .B(G92gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  AOI21_X1  g251(.A(new_n430_), .B1(new_n335_), .B2(new_n366_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n447_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n443_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n452_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n456_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT97), .B(new_n458_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n463_), .A2(KEYINPUT98), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT98), .B1(new_n463_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n429_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n452_), .A2(KEYINPUT32), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n448_), .A2(new_n456_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n422_), .A2(new_n410_), .A3(new_n423_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n425_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n470_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n445_), .A2(new_n447_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n390_), .A2(new_n391_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n454_), .B1(new_n476_), .B2(new_n453_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT32), .B(new_n452_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .A4(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n405_), .B1(new_n467_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT27), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n463_), .A2(new_n481_), .A3(new_n464_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n403_), .A2(new_n404_), .A3(new_n473_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n458_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT27), .A3(new_n457_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT102), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT102), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n482_), .A2(new_n483_), .A3(new_n488_), .A4(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n348_), .B1(new_n480_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n485_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n348_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n405_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n473_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .A4(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G29gat), .B(G36gat), .Z(new_n499_));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  INV_X1    g301(.A(G1gat), .ZN(new_n503_));
  INV_X1    g302(.A(G8gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G1gat), .B(G8gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n501_), .B(KEYINPUT15), .Z(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n501_), .A2(new_n508_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT79), .Z(new_n517_));
  NOR2_X1   g316(.A1(new_n511_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G113gat), .B(G141gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT80), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n522_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n296_), .B1(new_n498_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n526_), .ZN(new_n528_));
  AOI211_X1 g327(.A(KEYINPUT103), .B(new_n528_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n295_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n512_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT34), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n501_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n238_), .A2(new_n259_), .A3(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n531_), .A2(KEYINPUT73), .A3(new_n535_), .A4(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n534_), .B1(new_n531_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n512_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT69), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n543_), .B2(new_n263_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n545_));
  INV_X1    g344(.A(new_n537_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n538_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT74), .ZN(new_n550_));
  XOR2_X1   g349(.A(G134gat), .B(G162gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n552_), .A2(new_n553_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n548_), .A2(KEYINPUT75), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT75), .B1(new_n548_), .B2(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n560_));
  NAND2_X1  g359(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n548_), .A2(new_n556_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n548_), .A2(KEYINPUT75), .A3(new_n556_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n567_), .A2(KEYINPUT76), .A3(KEYINPUT37), .A4(new_n555_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n208_), .B(new_n508_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(KEYINPUT17), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n569_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n530_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n503_), .A3(new_n473_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n559_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n582_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n295_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n528_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n496_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(new_n587_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(G1324gat));
  AOI21_X1  g399(.A(new_n504_), .B1(new_n594_), .B2(new_n492_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT39), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n585_), .A2(new_n504_), .A3(new_n492_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n594_), .B2(new_n494_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n585_), .A2(new_n606_), .A3(new_n494_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1326gat));
  INV_X1    g409(.A(G22gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n594_), .B2(new_n405_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT42), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n585_), .A2(new_n611_), .A3(new_n405_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1327gat));
  NAND2_X1  g414(.A1(new_n589_), .A2(new_n582_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n295_), .B(new_n617_), .C1(new_n527_), .C2(new_n529_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n473_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n498_), .A2(new_n569_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT43), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n498_), .A2(new_n623_), .A3(new_n569_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n582_), .A3(new_n593_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n625_), .A2(KEYINPUT44), .A3(new_n582_), .A4(new_n593_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n473_), .A2(G29gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n620_), .B1(new_n630_), .B2(new_n631_), .ZN(G1328gat));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n492_), .A3(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n492_), .B(KEYINPUT105), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(G36gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n619_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT106), .B1(new_n618_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT45), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n634_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT46), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n634_), .B(KEYINPUT46), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1329gat));
  AOI21_X1  g447(.A(G43gat), .B1(new_n619_), .B2(new_n494_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n494_), .A2(G43gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n630_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT47), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1330gat));
  INV_X1    g453(.A(G50gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n619_), .A2(new_n655_), .A3(new_n405_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT107), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n630_), .A2(new_n405_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G50gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT107), .B(new_n655_), .C1(new_n630_), .C2(new_n405_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n295_), .A2(new_n526_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n498_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n583_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(G57gat), .A3(new_n496_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n590_), .A2(new_n591_), .A3(new_n662_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(new_n496_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(G57gat), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT108), .ZN(G1332gat));
  OAI21_X1  g468(.A(G64gat), .B1(new_n666_), .B2(new_n636_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT48), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n636_), .A2(G64gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n664_), .B2(new_n672_), .ZN(G1333gat));
  OAI21_X1  g472(.A(G71gat), .B1(new_n666_), .B2(new_n348_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT49), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n348_), .A2(G71gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n664_), .B2(new_n676_), .ZN(G1334gat));
  OAI21_X1  g476(.A(G78gat), .B1(new_n666_), .B2(new_n495_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT50), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n495_), .A2(G78gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n664_), .B2(new_n680_), .ZN(G1335gat));
  NAND2_X1  g480(.A1(new_n662_), .A2(new_n582_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n496_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n663_), .A2(new_n617_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n496_), .A2(G85gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(G1336gat));
  OAI21_X1  g487(.A(G92gat), .B1(new_n684_), .B2(new_n636_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n493_), .A2(G92gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n690_), .ZN(G1337gat));
  OAI21_X1  g490(.A(G99gat), .B1(new_n684_), .B2(new_n348_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n494_), .A2(new_n257_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n686_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g494(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n696_));
  INV_X1    g495(.A(new_n682_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n625_), .A2(new_n405_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n683_), .A2(new_n700_), .A3(new_n405_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n699_), .A2(G106gat), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT52), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n699_), .A2(new_n701_), .A3(new_n704_), .A4(G106gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n686_), .A2(G106gat), .A3(new_n495_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n696_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n696_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n707_), .B(new_n710_), .C1(new_n703_), .C2(new_n705_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1339gat));
  NAND2_X1  g511(.A1(new_n493_), .A2(new_n495_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n348_), .A3(new_n496_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT57), .ZN(new_n716_));
  INV_X1    g515(.A(new_n514_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n513_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(new_n522_), .C1(new_n717_), .C2(new_n518_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n720_), .A2(KEYINPUT114), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(KEYINPUT114), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n523_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n210_), .B1(new_n543_), .B2(new_n263_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n275_), .A3(new_n270_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n727_), .B2(KEYINPUT55), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT55), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n277_), .A2(KEYINPUT112), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(KEYINPUT55), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n265_), .A2(new_n266_), .A3(new_n276_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n278_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(KEYINPUT56), .A4(new_n285_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(new_n290_), .A3(new_n526_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n285_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT56), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n285_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(KEYINPUT113), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n724_), .B1(new_n737_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n716_), .B1(new_n743_), .B2(new_n589_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT115), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n716_), .C1(new_n743_), .C2(new_n589_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n737_), .A2(new_n742_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT57), .B(new_n559_), .C1(new_n749_), .C2(new_n724_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n723_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n285_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n285_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n569_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT58), .B(new_n751_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n569_), .B2(new_n756_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n750_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n582_), .B1(new_n748_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  INV_X1    g563(.A(new_n569_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n293_), .A2(new_n294_), .A3(new_n526_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n591_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(KEYINPUT54), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n583_), .A2(KEYINPUT111), .A3(new_n769_), .A4(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n715_), .B1(new_n763_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G113gat), .B1(new_n773_), .B2(new_n526_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n715_), .A2(KEYINPUT59), .ZN(new_n775_));
  INV_X1    g574(.A(new_n759_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n562_), .A2(new_n568_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n757_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n569_), .A2(new_n756_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT116), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n743_), .A2(new_n589_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n778_), .A2(new_n780_), .B1(KEYINPUT57), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n591_), .B1(new_n782_), .B2(new_n744_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n768_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n775_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n773_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n528_), .A2(KEYINPUT117), .ZN(new_n789_));
  MUX2_X1   g588(.A(KEYINPUT117), .B(new_n789_), .S(G113gat), .Z(new_n790_));
  AOI21_X1  g589(.A(new_n774_), .B1(new_n788_), .B2(new_n790_), .ZN(G1340gat));
  NOR2_X1   g590(.A1(new_n295_), .A2(KEYINPUT60), .ZN(new_n792_));
  MUX2_X1   g591(.A(new_n792_), .B(KEYINPUT60), .S(G120gat), .Z(new_n793_));
  AND2_X1   g592(.A1(new_n773_), .A2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT118), .Z(new_n795_));
  OAI21_X1  g594(.A(G120gat), .B1(new_n787_), .B2(new_n295_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1341gat));
  OAI211_X1 g596(.A(new_n591_), .B(new_n785_), .C1(new_n773_), .C2(new_n786_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G127gat), .ZN(new_n799_));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n773_), .A2(new_n800_), .A3(new_n591_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n804_), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1342gat));
  OAI21_X1  g605(.A(G134gat), .B1(new_n787_), .B2(new_n765_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n773_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n559_), .A2(G134gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(G1343gat));
  NAND2_X1  g609(.A1(new_n763_), .A2(new_n772_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n494_), .A2(new_n495_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n473_), .A3(new_n636_), .A4(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n528_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n372_), .ZN(G1344gat));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n295_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(new_n373_), .ZN(G1345gat));
  NOR2_X1   g616(.A1(new_n813_), .A2(new_n582_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT61), .B(G155gat), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n818_), .B(new_n819_), .Z(G1346gat));
  OAI21_X1  g619(.A(G162gat), .B1(new_n813_), .B2(new_n765_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n559_), .A2(G162gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n813_), .B2(new_n822_), .ZN(G1347gat));
  NOR3_X1   g622(.A1(new_n636_), .A2(new_n473_), .A3(new_n348_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n495_), .A3(new_n526_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n744_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n582_), .B1(new_n762_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n772_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G169gat), .B1(new_n828_), .B2(KEYINPUT120), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT121), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n829_), .A3(new_n834_), .A4(G169gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n835_), .A3(KEYINPUT62), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT121), .B(new_n837_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT22), .B(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n828_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n838_), .A3(new_n840_), .ZN(G1348gat));
  NOR2_X1   g640(.A1(new_n783_), .A2(new_n784_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n824_), .A2(new_n495_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G176gat), .B1(new_n844_), .B2(new_n592_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n763_), .A2(new_n772_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n846_), .A2(KEYINPUT122), .A3(new_n405_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT122), .B1(new_n846_), .B2(new_n405_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n824_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n295_), .A2(new_n309_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  AND3_X1   g650(.A1(new_n844_), .A2(new_n591_), .A3(new_n314_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n847_), .A2(new_n591_), .A3(new_n824_), .A4(new_n848_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n323_), .ZN(G1350gat));
  OR4_X1    g653(.A1(new_n559_), .A2(new_n842_), .A3(new_n432_), .A4(new_n843_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n324_), .B1(new_n844_), .B2(new_n569_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(G1351gat));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n812_), .A2(new_n496_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT124), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n636_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n811_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n811_), .A2(new_n860_), .A3(new_n863_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G197gat), .B1(new_n867_), .B2(new_n526_), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n351_), .B(new_n528_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1352gat));
  OAI211_X1 g669(.A(new_n867_), .B(new_n592_), .C1(KEYINPUT126), .C2(new_n352_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n352_), .A2(KEYINPUT126), .ZN(new_n872_));
  INV_X1    g671(.A(new_n866_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n864_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n874_), .B2(new_n295_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(G1353gat));
  NOR2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT127), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n582_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n867_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n878_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n881_), .B(new_n882_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1354gat));
  OAI21_X1  g683(.A(G218gat), .B1(new_n874_), .B2(new_n765_), .ZN(new_n885_));
  INV_X1    g684(.A(G218gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n867_), .A2(new_n886_), .A3(new_n589_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1355gat));
endmodule


