//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_;
  AND2_X1   g000(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(G78gat), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G78gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT65), .A2(G71gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n204_), .B(new_n210_), .C1(KEYINPUT11), .C2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n214_));
  INV_X1    g013(.A(G57gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(G64gat), .ZN(new_n216_));
  INV_X1    g015(.A(G64gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(G57gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n204_), .A4(new_n210_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(KEYINPUT11), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n213_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n213_), .B2(new_n221_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G85gat), .B(G92gat), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT9), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT6), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT8), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT6), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n235_), .A2(KEYINPUT6), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244_));
  INV_X1    g043(.A(G99gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n228_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n230_), .B(new_n239_), .C1(new_n243_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n247_), .B(new_n246_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n230_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n237_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n226_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G85gat), .B(G92gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n248_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n236_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n249_), .B(KEYINPUT67), .C1(new_n264_), .C2(new_n251_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n230_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n251_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT67), .B1(new_n269_), .B2(new_n249_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n237_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n213_), .A2(new_n221_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n222_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n213_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n260_), .B1(new_n226_), .B2(new_n255_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n257_), .A2(new_n272_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n261_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G120gat), .B(G148gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G176gat), .B(G204gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n261_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT69), .B1(new_n288_), .B2(new_n289_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT13), .B1(new_n292_), .B2(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G190gat), .B(G218gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G134gat), .B(G162gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT36), .Z(new_n305_));
  NAND2_X1  g104(.A1(G232gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT34), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT35), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G29gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G43gat), .B(G50gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n255_), .B2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(KEYINPUT15), .Z(new_n313_));
  INV_X1    g112(.A(new_n237_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n316_), .B2(new_n265_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n307_), .A2(KEYINPUT35), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT71), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n312_), .B(new_n320_), .C1(new_n313_), .C2(new_n317_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n305_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT74), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n304_), .A2(KEYINPUT36), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n329_), .A3(new_n324_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(new_n305_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT37), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n322_), .A2(new_n324_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n305_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n335_), .A2(new_n336_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G8gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT76), .ZN(new_n341_));
  INV_X1    g140(.A(G1gat), .ZN(new_n342_));
  INV_X1    g141(.A(G8gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT14), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT75), .B(KEYINPUT14), .C1(new_n342_), .C2(new_n343_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G15gat), .B(G22gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n341_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G231gat), .A3(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(G231gat), .ZN(new_n355_));
  INV_X1    g154(.A(G233gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n352_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n226_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT17), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n357_), .A3(new_n226_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G155gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G183gat), .B(G211gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(KEYINPUT78), .A3(new_n362_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n368_), .A2(KEYINPUT17), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n339_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n353_), .A2(new_n313_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n350_), .A2(new_n351_), .A3(new_n311_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G229gat), .A2(G233gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n353_), .A2(new_n311_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n379_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G141gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G169gat), .B(G197gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT79), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n385_), .A3(new_n391_), .A4(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n382_), .A2(new_n385_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n301_), .A2(new_n377_), .A3(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G197gat), .B(G204gat), .Z(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT21), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT21), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n401_), .A2(new_n404_), .A3(new_n402_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT24), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(G176gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n419_), .A2(new_n409_), .A3(new_n408_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT26), .B(G190gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT25), .B(G183gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n416_), .B(new_n420_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n419_), .A2(KEYINPUT89), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(KEYINPUT89), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n427_), .A2(new_n428_), .B1(new_n418_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n413_), .A2(new_n414_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n431_), .A2(KEYINPUT90), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT90), .B1(new_n431_), .B2(new_n432_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n407_), .A2(new_n426_), .A3(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n436_), .A2(KEYINPUT20), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n424_), .A2(new_n421_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT80), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(KEYINPUT80), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n420_), .A3(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n415_), .B(KEYINPUT81), .Z(new_n445_));
  NOR2_X1   g244(.A1(new_n431_), .A2(new_n432_), .ZN(new_n446_));
  AOI21_X1  g245(.A(G176gat), .B1(KEYINPUT82), .B2(KEYINPUT22), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(new_n417_), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n444_), .A2(new_n445_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n407_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n437_), .A2(new_n440_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT91), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n426_), .A2(new_n435_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n450_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(KEYINPUT20), .C1(new_n450_), .C2(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n439_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n437_), .A2(new_n458_), .A3(new_n440_), .A4(new_n451_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G8gat), .B(G36gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n453_), .A2(new_n467_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n437_), .A2(new_n451_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n439_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n439_), .B2(new_n456_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n472_), .B1(new_n475_), .B2(new_n465_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n469_), .A2(new_n471_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G141gat), .ZN(new_n479_));
  INV_X1    g278(.A(G148gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G141gat), .A2(G148gat), .ZN(new_n482_));
  INV_X1    g281(.A(G155gat), .ZN(new_n483_));
  INV_X1    g282(.A(G162gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT1), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(G155gat), .B2(G162gat), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT1), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n481_), .B(new_n482_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G155gat), .B(G162gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n481_), .B1(new_n492_), .B2(KEYINPUT3), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n494_), .A2(new_n479_), .A3(new_n480_), .A4(KEYINPUT85), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  AND4_X1   g297(.A1(new_n493_), .A2(new_n495_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n488_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n500_));
  OR3_X1    g299(.A1(new_n500_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT28), .B1(new_n500_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n407_), .B1(KEYINPUT29), .B2(new_n500_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(G228gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(G228gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n356_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G78gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n228_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G22gat), .B(G50gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n505_), .A2(new_n506_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n478_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(G127gat), .B(G134gat), .Z(new_n521_));
  XOR2_X1   g320(.A(G113gat), .B(G120gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n523_), .B(new_n488_), .C1(new_n499_), .C2(new_n491_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n500_), .A2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT4), .B(new_n524_), .C1(new_n526_), .C2(KEYINPUT93), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n500_), .A2(new_n525_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n520_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n526_), .A2(new_n524_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n520_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G85gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT0), .B(G57gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n531_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n449_), .B(KEYINPUT30), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT83), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546_));
  INV_X1    g345(.A(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(G15gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n548_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(new_n544_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n523_), .B(KEYINPUT31), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n519_), .A2(new_n542_), .A3(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n466_), .A2(new_n468_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n540_), .A2(KEYINPUT33), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(new_n538_), .C1(new_n531_), .C2(new_n534_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n527_), .A2(new_n520_), .A3(new_n530_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT94), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n538_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n563_), .A2(KEYINPUT95), .A3(new_n567_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n571_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n469_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n475_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(KEYINPUT96), .Z(new_n578_));
  OAI211_X1 g377(.A(new_n541_), .B(new_n577_), .C1(new_n460_), .C2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n517_), .A2(new_n541_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n580_), .A2(new_n517_), .B1(new_n581_), .B2(new_n477_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n559_), .A2(KEYINPUT84), .A3(new_n560_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT84), .B1(new_n559_), .B2(new_n560_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n562_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n398_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT98), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n541_), .B(KEYINPUT99), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(G1gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT100), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n328_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n587_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n297_), .A2(new_n298_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n397_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n374_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n542_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n593_), .A2(KEYINPUT38), .A3(new_n595_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n598_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NAND4_X1  g406(.A1(new_n586_), .A2(new_n603_), .A3(new_n478_), .A4(new_n335_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(G8gat), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT102), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n610_), .A2(new_n615_), .A3(G8gat), .A4(new_n611_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(KEYINPUT39), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n589_), .A2(new_n343_), .A3(new_n478_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(KEYINPUT40), .A3(new_n617_), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1325gat));
  INV_X1    g422(.A(G15gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n589_), .A2(new_n624_), .A3(new_n585_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(new_n585_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G15gat), .B1(new_n604_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n626_), .A2(new_n629_), .A3(new_n630_), .A4(new_n631_), .ZN(G1326gat));
  NAND3_X1  g431(.A1(new_n600_), .A2(new_n518_), .A3(new_n603_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G22gat), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT104), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT104), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT42), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n589_), .A2(new_n638_), .A3(new_n518_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT42), .B1(new_n635_), .B2(new_n636_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  NOR2_X1   g441(.A1(new_n375_), .A2(new_n335_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT108), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n602_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n586_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(G29gat), .A3(new_n542_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n602_), .A2(new_n375_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n332_), .A2(new_n338_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n599_), .B2(KEYINPUT37), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT43), .B1(new_n339_), .B2(KEYINPUT105), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n586_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n586_), .B2(new_n650_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  INV_X1    g456(.A(new_n590_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n648_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .A4(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(G29gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT106), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT107), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  AND4_X1   g463(.A1(KEYINPUT107), .A2(new_n663_), .A3(G29gat), .A4(new_n660_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n647_), .B1(new_n664_), .B2(new_n665_), .ZN(G1328gat));
  NAND3_X1  g465(.A1(new_n656_), .A2(new_n478_), .A3(new_n659_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n477_), .A2(G36gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n645_), .A2(new_n586_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT45), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT109), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT109), .B(new_n674_), .C1(new_n668_), .C2(new_n671_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1329gat));
  NAND4_X1  g475(.A1(new_n656_), .A2(G43gat), .A3(new_n561_), .A4(new_n659_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n547_), .B1(new_n646_), .B2(new_n627_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g479(.A1(new_n656_), .A2(G50gat), .A3(new_n518_), .A4(new_n659_), .ZN(new_n681_));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n646_), .B2(new_n517_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1331gat));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n301_), .A2(new_n374_), .A3(new_n397_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n600_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n586_), .A3(new_n335_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT111), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n687_), .A2(new_n541_), .A3(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n587_), .A2(new_n397_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT110), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n376_), .A2(new_n601_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n658_), .A2(new_n215_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n215_), .A2(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(G1332gat));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n478_), .A3(new_n687_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G64gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G64gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n478_), .A2(new_n217_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n699_), .A2(new_n700_), .B1(new_n694_), .B2(new_n701_), .ZN(G1333gat));
  NAND3_X1  g501(.A1(new_n689_), .A2(new_n585_), .A3(new_n687_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G71gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G71gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n585_), .A2(new_n206_), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n705_), .A2(new_n706_), .B1(new_n694_), .B2(new_n707_), .ZN(G1334gat));
  NAND4_X1  g507(.A1(new_n692_), .A2(new_n208_), .A3(new_n518_), .A4(new_n693_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n689_), .A2(new_n518_), .A3(new_n687_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G78gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G78gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n709_), .B(KEYINPUT112), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n601_), .A2(new_n375_), .A3(new_n397_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n542_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n644_), .A2(new_n301_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n692_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n658_), .A2(new_n232_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1336gat));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n692_), .A2(new_n478_), .A3(new_n722_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n728_), .B2(G92gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(KEYINPUT113), .A3(new_n233_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n720_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n477_), .A2(new_n233_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n729_), .A2(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(G1337gat));
  NAND4_X1  g532(.A1(new_n692_), .A2(new_n561_), .A3(new_n227_), .A4(new_n722_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n585_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n245_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g537(.A1(new_n518_), .A2(new_n228_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n518_), .B(new_n719_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n723_), .A2(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g544(.A(G113gat), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT59), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n372_), .A2(new_n397_), .A3(new_n373_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n749_), .A2(new_n297_), .A3(KEYINPUT114), .A4(new_n298_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n748_), .B1(new_n754_), .B2(new_n339_), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT54), .B(new_n650_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT55), .A4(new_n279_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT115), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n271_), .A2(new_n276_), .B1(new_n257_), .B2(new_n272_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT55), .A4(new_n278_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n277_), .A2(new_n256_), .A3(new_n279_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n765_), .A2(new_n280_), .B1(new_n766_), .B2(new_n260_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(KEYINPUT116), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n287_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT116), .B1(new_n764_), .B2(new_n767_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n758_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n764_), .A2(new_n767_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n287_), .A4(new_n768_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT118), .B(new_n758_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n378_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n381_), .B1(new_n384_), .B2(new_n379_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n395_), .A3(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n393_), .A2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n289_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n650_), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n293_), .A2(new_n783_), .A3(new_n295_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n397_), .A2(new_n289_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n771_), .B2(new_n777_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT117), .B(new_n791_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n335_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n335_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n789_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n757_), .B1(new_n800_), .B2(new_n374_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n519_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n561_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n802_), .A2(new_n590_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n747_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n339_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n807_), .A2(new_n788_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n375_), .B1(new_n808_), .B2(new_n799_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT59), .B(new_n804_), .C1(new_n809_), .C2(new_n757_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n746_), .B1(new_n811_), .B2(new_n397_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n801_), .A2(new_n805_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n397_), .A2(new_n746_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT119), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  INV_X1    g617(.A(new_n397_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n820_));
  OAI221_X1 g619(.A(new_n818_), .B1(new_n814_), .B2(new_n815_), .C1(new_n820_), .C2(new_n746_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n813_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n301_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  OAI21_X1  g626(.A(G120gat), .B1(new_n826_), .B2(KEYINPUT120), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n811_), .B2(new_n375_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n375_), .A2(new_n830_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n814_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT121), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n374_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n836_));
  OAI221_X1 g635(.A(new_n835_), .B1(new_n814_), .B2(new_n832_), .C1(new_n836_), .C2(new_n830_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n813_), .B2(new_n599_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT122), .B(G134gat), .Z(new_n840_));
  NOR2_X1   g639(.A1(new_n339_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n811_), .B2(new_n841_), .ZN(G1343gat));
  NOR4_X1   g641(.A1(new_n585_), .A2(new_n517_), .A3(new_n478_), .A4(new_n590_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n801_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n397_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT124), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n848_), .A3(new_n397_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT123), .B(G141gat), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1344gat));
  INV_X1    g652(.A(new_n845_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n301_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n480_), .ZN(G1345gat));
  NAND2_X1  g655(.A1(new_n845_), .A2(new_n375_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  OAI21_X1  g658(.A(G162gat), .B1(new_n854_), .B2(new_n339_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n845_), .A2(new_n484_), .A3(new_n599_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1347gat));
  NOR2_X1   g661(.A1(new_n801_), .A2(new_n477_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n627_), .A2(new_n518_), .A3(new_n658_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n397_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(G169gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(G169gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n864_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n397_), .A2(new_n429_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT125), .Z(new_n871_));
  OAI22_X1  g670(.A1(new_n867_), .A2(new_n868_), .B1(new_n869_), .B2(new_n871_), .ZN(G1348gat));
  OAI21_X1  g671(.A(G176gat), .B1(new_n869_), .B2(new_n301_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n299_), .A2(new_n418_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n869_), .B2(new_n874_), .ZN(G1349gat));
  NAND3_X1  g674(.A1(new_n863_), .A2(new_n375_), .A3(new_n864_), .ZN(new_n876_));
  MUX2_X1   g675(.A(new_n424_), .B(G183gat), .S(new_n876_), .Z(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n869_), .B2(new_n339_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n335_), .A2(new_n423_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n869_), .B2(new_n879_), .ZN(G1351gat));
  NAND3_X1  g679(.A1(new_n863_), .A2(new_n581_), .A3(new_n627_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n819_), .ZN(new_n882_));
  INV_X1    g681(.A(G197gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1352gat));
  NOR2_X1   g683(.A1(new_n881_), .A2(new_n301_), .ZN(new_n885_));
  INV_X1    g684(.A(G204gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1353gat));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n888_));
  INV_X1    g687(.A(G211gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n375_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n881_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n889_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT126), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n891_), .B(new_n893_), .ZN(G1354gat));
  OAI21_X1  g693(.A(G218gat), .B1(new_n881_), .B2(new_n339_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n335_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n881_), .B2(new_n896_), .ZN(G1355gat));
endmodule


