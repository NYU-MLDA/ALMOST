//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n207_), .A3(new_n210_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT66), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT66), .B1(new_n212_), .B2(new_n214_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n221_), .B(new_n206_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n206_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n224_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n220_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n231_), .B2(new_n203_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n215_), .A3(new_n228_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n202_), .A2(KEYINPUT8), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n216_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(G71gat), .A2(G78gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G71gat), .A2(G78gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G57gat), .B(G64gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT11), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n244_), .B2(KEYINPUT11), .ZN(new_n247_));
  INV_X1    g046(.A(G64gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G57gat), .ZN(new_n249_));
  INV_X1    g048(.A(G57gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G64gat), .ZN(new_n251_));
  AND4_X1   g050(.A1(new_n246_), .A2(new_n249_), .A3(new_n251_), .A4(KEYINPUT11), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n245_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n251_), .A3(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT68), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n251_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n249_), .A2(new_n251_), .A3(new_n246_), .A4(KEYINPUT11), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n243_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n240_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n253_), .A2(new_n260_), .A3(KEYINPUT69), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n234_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n236_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n227_), .B1(new_n226_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n223_), .B1(new_n221_), .B2(new_n206_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT67), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n224_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n202_), .B1(new_n276_), .B2(new_n220_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n270_), .B1(new_n277_), .B2(new_n217_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n268_), .B1(new_n278_), .B2(new_n216_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n279_), .B2(KEYINPUT12), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n216_), .A3(new_n268_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G230gat), .A2(G233gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(KEYINPUT70), .A3(new_n282_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n280_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n268_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n240_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n289_), .B2(new_n281_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G120gat), .B(G148gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G176gat), .B(G204gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n291_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT13), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(G29gat), .B(G36gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT74), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(KEYINPUT74), .ZN(new_n315_));
  XOR2_X1   g114(.A(G43gat), .B(G50gat), .Z(new_n316_));
  OR3_X1    g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n312_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G229gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n319_), .B(KEYINPUT15), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n310_), .B(new_n311_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n312_), .A2(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n321_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n303_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n328_), .A2(new_n326_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n335_), .A2(KEYINPUT81), .A3(new_n323_), .A4(new_n332_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n332_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(KEYINPUT80), .A3(new_n323_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n334_), .A2(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G127gat), .B(G155gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(G183gat), .B(G211gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G231gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n325_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n261_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n352_), .B2(KEYINPUT69), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(KEYINPUT69), .B2(new_n352_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n352_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n346_), .A2(new_n347_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n302_), .A2(new_n341_), .A3(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n363_), .A2(KEYINPUT99), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(KEYINPUT99), .ZN(new_n365_));
  XOR2_X1   g164(.A(G211gat), .B(G218gat), .Z(new_n366_));
  INV_X1    g165(.A(G197gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G204gat), .ZN(new_n368_));
  INV_X1    g167(.A(G204gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G197gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n366_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n367_), .A3(G204gat), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT21), .B(new_n376_), .C1(new_n371_), .C2(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n372_), .A2(new_n373_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n374_), .A2(new_n377_), .B1(new_n378_), .B2(new_n366_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT88), .B1(new_n391_), .B2(KEYINPUT1), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n392_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(KEYINPUT1), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT87), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n391_), .A2(new_n401_), .A3(KEYINPUT1), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n386_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n384_), .B(KEYINPUT3), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n382_), .B(KEYINPUT2), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n407_), .A2(new_n391_), .A3(new_n397_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n381_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT93), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n379_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n410_), .B2(new_n409_), .ZN(new_n412_));
  INV_X1    g211(.A(G233gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n379_), .A2(new_n417_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n400_), .A2(new_n402_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n392_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n385_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n408_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT89), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n419_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G22gat), .B(G50gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT28), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n427_), .A2(new_n433_), .A3(new_n428_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n436_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n440_), .B2(new_n434_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n431_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n418_), .A2(new_n429_), .A3(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n432_), .A2(new_n439_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n439_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n418_), .A2(new_n429_), .A3(new_n442_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n418_), .B2(new_n429_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT24), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(G169gat), .B2(G176gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453_));
  INV_X1    g252(.A(G169gat), .ZN(new_n454_));
  INV_X1    g253(.A(G176gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT83), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT25), .B(G183gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT26), .B(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT23), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT23), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n459_), .A2(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n451_), .A2(new_n456_), .A3(new_n466_), .A4(new_n452_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n456_), .A2(new_n452_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n450_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n458_), .A2(new_n465_), .A3(new_n467_), .A4(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n463_), .B2(new_n461_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n463_), .B2(new_n461_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT22), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n455_), .B1(new_n474_), .B2(KEYINPUT84), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(G169gat), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n475_), .A2(G169gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n479_), .B(KEYINPUT30), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT85), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(KEYINPUT85), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G43gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G15gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  MUX2_X1   g286(.A(new_n481_), .B(new_n482_), .S(new_n487_), .Z(new_n488_));
  XNOR2_X1  g287(.A(G127gat), .B(G134gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G113gat), .B(G120gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT31), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n488_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT22), .B(G169gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n455_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n473_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n462_), .A2(new_n464_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n454_), .A2(new_n455_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(KEYINPUT24), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT94), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n499_), .B(new_n503_), .C1(KEYINPUT24), .C2(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n459_), .A2(new_n460_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n506_), .A2(new_n457_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n498_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n494_), .B1(new_n508_), .B2(new_n379_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT19), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n374_), .A2(new_n377_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n378_), .A2(new_n366_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n479_), .B2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n479_), .A2(new_n516_), .A3(new_n513_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n509_), .B(new_n512_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G8gat), .B(G36gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT18), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n379_), .A2(new_n470_), .A3(new_n478_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n524_), .B(KEYINPUT20), .C1(new_n508_), .C2(new_n379_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n511_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n519_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n525_), .A2(new_n511_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n509_), .B1(new_n518_), .B2(new_n517_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n511_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(new_n523_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT98), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n532_), .A2(new_n535_), .A3(new_n523_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n529_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n523_), .B1(new_n519_), .B2(new_n526_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n527_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n424_), .A2(new_n426_), .A3(new_n491_), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n404_), .A2(new_n408_), .A3(new_n491_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n541_), .A2(KEYINPUT4), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n424_), .A2(new_n426_), .A3(new_n544_), .A4(new_n491_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G225gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT96), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n541_), .A2(KEYINPUT97), .A3(new_n542_), .A4(new_n546_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n541_), .A2(KEYINPUT4), .A3(new_n542_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n547_), .A4(new_n545_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G29gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G85gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT0), .B(G57gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n549_), .A2(new_n554_), .A3(new_n562_), .A4(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR4_X1   g365(.A1(new_n449_), .A2(new_n493_), .A3(new_n540_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n540_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n449_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n523_), .A2(KEYINPUT32), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n519_), .A2(new_n571_), .A3(new_n526_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n532_), .B2(new_n571_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n555_), .A2(new_n546_), .A3(new_n545_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n541_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n563_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n527_), .A2(new_n538_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n565_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n549_), .A2(new_n557_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(KEYINPUT33), .A3(new_n562_), .A4(new_n554_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n566_), .A2(new_n574_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n570_), .B1(new_n584_), .B2(new_n449_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n567_), .B1(new_n585_), .B2(new_n493_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n324_), .A2(new_n240_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n278_), .A2(new_n319_), .A3(new_n216_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n594_), .A2(new_n595_), .B1(KEYINPUT36), .B2(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT35), .ZN(new_n599_));
  XOR2_X1   g398(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(KEYINPUT75), .A3(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n597_), .B2(KEYINPUT75), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n591_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n596_), .A2(new_n602_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n607_), .A2(new_n590_), .A3(new_n604_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n364_), .A2(new_n365_), .A3(new_n586_), .A4(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT100), .Z(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n569_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n302_), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n606_), .A2(new_n608_), .B1(KEYINPUT76), .B2(KEYINPUT37), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n603_), .A2(new_n591_), .A3(new_n605_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n590_), .B1(new_n607_), .B2(new_n604_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n362_), .ZN(new_n621_));
  NOR4_X1   g420(.A1(new_n586_), .A2(new_n340_), .A3(new_n613_), .A4(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n304_), .A3(new_n566_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n612_), .A2(new_n624_), .ZN(G1324gat));
  AOI21_X1  g424(.A(new_n305_), .B1(new_n610_), .B2(new_n540_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT39), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n305_), .A3(new_n540_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n611_), .B2(new_n493_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(G15gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n493_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n622_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(G1326gat));
  NAND2_X1  g437(.A1(new_n444_), .A2(new_n448_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G22gat), .B1(new_n611_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT42), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(G22gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT101), .Z(new_n643_));
  NAND2_X1  g442(.A1(new_n622_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n609_), .A2(new_n361_), .ZN(new_n647_));
  NOR4_X1   g446(.A1(new_n586_), .A2(new_n340_), .A3(new_n613_), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n566_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n302_), .A2(new_n341_), .A3(new_n361_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n620_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n566_), .A2(new_n574_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n581_), .A2(new_n583_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n639_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n636_), .B1(new_n657_), .B2(new_n570_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n658_), .B2(new_n567_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT43), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n449_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n540_), .A2(new_n639_), .A3(new_n566_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n493_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n449_), .A2(new_n540_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n569_), .A3(new_n636_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n620_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(KEYINPUT102), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n652_), .B1(new_n661_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT103), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n667_), .B2(KEYINPUT102), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n660_), .B(KEYINPUT43), .C1(new_n586_), .C2(new_n620_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n651_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n672_), .A2(new_n677_), .B1(KEYINPUT44), .B2(new_n676_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n566_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n646_), .B(new_n650_), .C1(new_n679_), .C2(new_n649_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n649_), .B1(new_n678_), .B2(new_n566_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n650_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT104), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n648_), .A2(new_n685_), .A3(new_n540_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT45), .Z(new_n687_));
  AOI21_X1  g486(.A(new_n568_), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT103), .B1(new_n670_), .B2(new_n671_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n676_), .A2(new_n673_), .A3(KEYINPUT44), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n691_), .B2(G36gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n692_), .A2(KEYINPUT105), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n652_), .C1(new_n661_), .C2(new_n669_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n540_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n677_), .B2(new_n672_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n685_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n693_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n695_), .A2(new_n702_), .ZN(G1329gat));
  AOI21_X1  g502(.A(G43gat), .B1(new_n648_), .B2(new_n636_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n636_), .A2(G43gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n678_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n648_), .B2(new_n449_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n449_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n678_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(G1331gat));
  NAND3_X1  g512(.A1(new_n613_), .A2(new_n340_), .A3(new_n362_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n586_), .A2(new_n714_), .A3(new_n609_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(G57gat), .A3(new_n566_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n586_), .A2(new_n341_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n621_), .A2(new_n302_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n250_), .B1(new_n720_), .B2(new_n569_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT109), .Z(G1332gat));
  AOI21_X1  g523(.A(new_n248_), .B1(new_n715_), .B2(new_n540_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n540_), .A2(new_n248_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT111), .Z(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n720_), .B2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n715_), .B2(new_n636_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  INV_X1    g532(.A(new_n720_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n731_), .A3(new_n636_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT112), .Z(G1334gat));
  INV_X1    g536(.A(G78gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n715_), .B2(new_n449_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n738_), .A3(new_n449_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NOR4_X1   g541(.A1(new_n586_), .A2(new_n341_), .A3(new_n302_), .A4(new_n647_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n566_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT113), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n613_), .A2(new_n340_), .A3(new_n361_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n569_), .A2(new_n208_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n743_), .A2(new_n209_), .A3(new_n540_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n747_), .A2(new_n540_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n209_), .ZN(G1337gat));
  AND3_X1   g551(.A1(new_n743_), .A2(new_n636_), .A3(new_n205_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n221_), .B1(new_n747_), .B2(new_n636_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n753_), .B(new_n754_), .C1(KEYINPUT114), .C2(KEYINPUT51), .ZN(new_n755_));
  NOR2_X1   g554(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1338gat));
  AOI21_X1  g556(.A(new_n206_), .B1(new_n747_), .B2(new_n449_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n758_), .A2(KEYINPUT52), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n743_), .A2(new_n206_), .A3(new_n449_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT115), .Z(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(KEYINPUT52), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g563(.A1(new_n302_), .A2(new_n340_), .A3(new_n362_), .A4(new_n620_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n332_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n327_), .A2(new_n322_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n326_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n296_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n287_), .A2(new_n290_), .A3(new_n773_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n772_), .B(new_n774_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT55), .B1(new_n287_), .B2(KEYINPUT116), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n289_), .A2(new_n262_), .B1(new_n240_), .B2(new_n263_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n286_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT70), .B1(new_n281_), .B2(new_n282_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n281_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(G230gat), .A3(G233gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n773_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n773_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n775_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n620_), .B1(new_n768_), .B2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n787_), .A2(new_n788_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n775_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n789_), .B2(new_n768_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n340_), .A2(new_n774_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n772_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n298_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n609_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT117), .B(new_n609_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n795_), .B(new_n801_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n767_), .B1(new_n806_), .B2(new_n361_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n665_), .A2(new_n566_), .A3(new_n636_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n341_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT59), .B1(new_n807_), .B2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n795_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT119), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n795_), .B(new_n815_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n801_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n767_), .B1(new_n817_), .B2(new_n361_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n808_), .A2(KEYINPUT59), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n811_), .B(new_n812_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n801_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n813_), .B2(KEYINPUT119), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n362_), .B1(new_n824_), .B2(new_n816_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n819_), .B1(new_n825_), .B2(new_n767_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n811_), .B1(new_n826_), .B2(new_n812_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n822_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n340_), .A2(KEYINPUT121), .ZN(new_n829_));
  MUX2_X1   g628(.A(KEYINPUT121), .B(new_n829_), .S(G113gat), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n810_), .B1(new_n828_), .B2(new_n830_), .ZN(G1340gat));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n302_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n809_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n832_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n826_), .A2(new_n613_), .A3(new_n812_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n809_), .A2(new_n838_), .A3(new_n362_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n822_), .A2(new_n827_), .A3(new_n361_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n809_), .A2(new_n842_), .A3(new_n609_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n822_), .A2(new_n827_), .A3(new_n620_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n807_), .A2(new_n636_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n569_), .A2(new_n540_), .A3(new_n639_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n341_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n613_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g651(.A1(new_n846_), .A2(new_n362_), .A3(new_n847_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n848_), .A2(new_n860_), .A3(new_n609_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n848_), .A2(new_n653_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1347gat));
  INV_X1    g662(.A(new_n818_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n568_), .A2(new_n449_), .A3(new_n493_), .A4(new_n566_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n496_), .A3(new_n341_), .A4(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n454_), .A2(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n341_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n818_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n341_), .B(new_n865_), .C1(new_n825_), .C2(new_n767_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT123), .A3(new_n867_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n872_), .B2(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n871_), .B(new_n873_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT124), .B(new_n874_), .C1(new_n872_), .C2(G169gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n866_), .B1(new_n877_), .B2(new_n878_), .ZN(G1348gat));
  INV_X1    g678(.A(new_n767_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n806_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n362_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(new_n865_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(G176gat), .A3(new_n613_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n864_), .A2(new_n865_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G176gat), .B1(new_n887_), .B2(new_n613_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1349gat));
  AOI21_X1  g688(.A(G183gat), .B1(new_n883_), .B2(new_n362_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n361_), .A2(new_n459_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n887_), .B2(new_n891_), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n887_), .A2(new_n653_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G190gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n887_), .A2(new_n460_), .A3(new_n609_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n568_), .A2(new_n566_), .A3(new_n639_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n882_), .A2(new_n493_), .A3(new_n897_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n900_));
  OAI211_X1 g699(.A(G197gat), .B(new_n341_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n898_), .B(KEYINPUT126), .ZN(new_n903_));
  AOI21_X1  g702(.A(G197gat), .B1(new_n903_), .B2(new_n341_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n613_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G204gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n903_), .A2(new_n369_), .A3(new_n613_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1353gat));
  AOI21_X1  g708(.A(new_n361_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT127), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n903_), .A2(new_n913_), .A3(new_n910_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n903_), .A2(new_n918_), .A3(new_n609_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n903_), .A2(new_n653_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n918_), .ZN(G1355gat));
endmodule


