//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n205_), .A3(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n206_), .A2(KEYINPUT25), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G183gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(new_n212_), .B2(new_n213_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G176gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(KEYINPUT24), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n215_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT79), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(new_n215_), .C1(new_n226_), .C2(new_n229_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n234_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n245_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G15gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT30), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n255_), .B(new_n258_), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n240_), .A2(new_n241_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G155gat), .B(G162gat), .Z(new_n263_));
  INV_X1    g062(.A(G141gat), .ZN(new_n264_));
  INV_X1    g063(.A(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT3), .B1(new_n266_), .B2(KEYINPUT83), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT2), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n266_), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n263_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n245_), .A2(new_n246_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n255_), .B2(new_n279_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT93), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n244_), .B1(new_n253_), .B2(new_n249_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n250_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n279_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n281_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT92), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n282_), .A2(new_n292_), .A3(KEYINPUT4), .ZN(new_n293_));
  INV_X1    g092(.A(new_n288_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n285_), .B1(new_n297_), .B2(new_n284_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G85gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G57gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n284_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n290_), .A2(KEYINPUT92), .B1(new_n294_), .B2(new_n295_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n293_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n307_), .A2(new_n302_), .A3(new_n285_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n211_), .A2(G169gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n213_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT89), .B1(new_n212_), .B2(new_n213_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G169gat), .A3(G176gat), .ZN(new_n317_));
  AND4_X1   g116(.A1(new_n209_), .A2(new_n314_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT88), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT24), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n225_), .B(new_n324_), .C1(new_n228_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n219_), .A2(new_n221_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n219_), .A2(new_n221_), .A3(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n216_), .A2(new_n218_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n318_), .B1(new_n327_), .B2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(KEYINPUT21), .A3(new_n336_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT90), .B1(new_n334_), .B2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n209_), .A2(new_n314_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n326_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT90), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n344_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n231_), .A2(new_n345_), .A3(new_n233_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT20), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n353_), .B2(KEYINPUT20), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n311_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n234_), .A2(new_n345_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n349_), .B2(new_n344_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n359_), .A2(new_n311_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT18), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n358_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT91), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT91), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n358_), .A2(new_n361_), .A3(new_n371_), .A4(new_n366_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT96), .B(KEYINPUT27), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT84), .B(KEYINPUT29), .Z(new_n375_));
  AOI21_X1  g174(.A(new_n345_), .B1(new_n279_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n377_), .A3(new_n344_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT85), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n385_));
  XOR2_X1   g184(.A(G22gat), .B(G50gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT28), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n385_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n381_), .A2(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n383_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n384_), .A2(new_n390_), .A3(new_n383_), .A4(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n311_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT95), .B(new_n311_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n357_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n397_), .B(new_n398_), .C1(new_n311_), .C2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n367_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n309_), .A2(new_n374_), .A3(new_n394_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n262_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n370_), .A2(new_n372_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT33), .B(new_n302_), .C1(new_n307_), .C2(new_n285_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n302_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n297_), .B2(new_n284_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n358_), .A2(new_n361_), .A3(new_n414_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n401_), .A2(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI221_X1 g217(.A(new_n418_), .B1(new_n417_), .B2(new_n416_), .C1(new_n304_), .C2(new_n308_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n394_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n404_), .A2(new_n405_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n406_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n374_), .A2(new_n403_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n374_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n394_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT99), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n262_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n374_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT98), .B1(new_n374_), .B2(new_n403_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n421_), .B(new_n431_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT99), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n424_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT72), .B(G15gat), .ZN(new_n438_));
  INV_X1    g237(.A(G22gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT73), .B(G8gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT14), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G8gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G29gat), .B(G36gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT70), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G43gat), .B(G50gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n451_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT15), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n451_), .B(new_n452_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT15), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n449_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G229gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n447_), .A2(new_n448_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n449_), .A2(new_n454_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n457_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT76), .B1(new_n467_), .B2(new_n461_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n469_), .B(new_n460_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G169gat), .B(G197gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n464_), .B(new_n474_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT77), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n479_), .A3(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT78), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n437_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G230gat), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(G85gat), .B2(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT9), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT64), .B(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n493_), .B2(KEYINPUT65), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(KEYINPUT65), .B2(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT10), .B(G99gat), .Z(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  NOR2_X1   g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n503_), .B1(new_n506_), .B2(new_n498_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT8), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n502_), .A2(new_n508_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n487_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT66), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n521_), .B(new_n487_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n502_), .A2(new_n508_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n515_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(KEYINPUT12), .A3(new_n516_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n518_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n487_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OR3_X1    g329(.A1(new_n523_), .A2(KEYINPUT69), .A3(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G120gat), .B(G148gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT67), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT69), .B1(new_n523_), .B2(new_n530_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n531_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n485_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n515_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n462_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G127gat), .B(G155gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT17), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT75), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n551_), .A2(new_n559_), .A3(new_n555_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n456_), .A2(new_n458_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n502_), .A2(new_n508_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT34), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n524_), .A2(new_n454_), .B1(KEYINPUT35), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT35), .B(new_n566_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(KEYINPUT36), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n578_), .B(KEYINPUT37), .C1(new_n573_), .C2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(KEYINPUT71), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n572_), .B2(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n581_), .A2(new_n583_), .B1(new_n577_), .B2(new_n573_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n584_), .B2(KEYINPUT37), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n547_), .A2(new_n561_), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n484_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n309_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n442_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT38), .ZN(new_n590_));
  INV_X1    g389(.A(new_n481_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n546_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n561_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n546_), .A2(KEYINPUT100), .A3(new_n591_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n584_), .B(KEYINPUT101), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n597_), .A2(new_n437_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n442_), .B1(new_n600_), .B2(new_n588_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n590_), .B1(new_n603_), .B2(new_n604_), .ZN(G1324gat));
  XNOR2_X1  g404(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n437_), .A2(new_n599_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n427_), .A2(new_n428_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612_));
  OAI21_X1  g411(.A(G8gat), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT103), .B1(new_n600_), .B2(new_n609_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT39), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n612_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n600_), .A2(KEYINPUT103), .A3(new_n609_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .A4(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n587_), .A2(new_n609_), .A3(new_n441_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n606_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n606_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n621_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n623_), .B(new_n624_), .C1(new_n615_), .C2(new_n619_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n262_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n587_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT105), .ZN(new_n630_));
  INV_X1    g429(.A(new_n600_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n631_), .B2(new_n262_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(new_n633_), .A3(new_n634_), .ZN(G1326gat));
  XNOR2_X1  g434(.A(new_n394_), .B(KEYINPUT106), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n587_), .A2(new_n439_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n439_), .B1(new_n600_), .B2(new_n636_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT42), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  NAND2_X1  g441(.A1(new_n584_), .A2(new_n561_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n547_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n484_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G29gat), .A3(new_n309_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n594_), .A2(new_n561_), .A3(new_n596_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n404_), .A2(new_n405_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n394_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n404_), .A2(new_n405_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n650_), .B(new_n262_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n430_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n435_), .A2(KEYINPUT99), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n585_), .B(KEYINPUT107), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n649_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n585_), .A2(new_n649_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n432_), .A2(new_n436_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n653_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n648_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n648_), .C1(new_n658_), .C2(new_n661_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n588_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n646_), .B1(new_n666_), .B2(G29gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT108), .ZN(G1328gat));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n585_), .B(KEYINPUT107), .Z(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n437_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n661_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n674_), .B2(new_n648_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n665_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n670_), .B1(new_n677_), .B2(new_n609_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n484_), .A2(new_n670_), .A3(new_n609_), .A4(new_n644_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT45), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n669_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n675_), .A2(new_n676_), .A3(new_n608_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n680_), .B(KEYINPUT46), .C1(new_n683_), .C2(new_n670_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1329gat));
  NOR2_X1   g484(.A1(new_n262_), .A2(new_n236_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n664_), .A2(new_n665_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT109), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n664_), .A2(new_n689_), .A3(new_n665_), .A4(new_n686_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n236_), .B1(new_n645_), .B2(new_n262_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n688_), .A2(new_n694_), .A3(new_n690_), .A4(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  NOR3_X1   g495(.A1(new_n675_), .A2(new_n676_), .A3(new_n421_), .ZN(new_n697_));
  INV_X1    g496(.A(G50gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n636_), .A2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT110), .Z(new_n700_));
  OAI22_X1  g499(.A1(new_n697_), .A2(new_n698_), .B1(new_n645_), .B2(new_n700_), .ZN(G1331gat));
  NAND3_X1  g500(.A1(new_n656_), .A2(new_n481_), .A3(new_n547_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n561_), .A3(new_n585_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n588_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n546_), .A2(new_n482_), .A3(new_n561_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n607_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n309_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n708_), .B2(new_n609_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n704_), .A2(new_n712_), .A3(new_n609_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n708_), .B2(new_n628_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT49), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n704_), .A2(new_n717_), .A3(new_n628_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n708_), .B2(new_n636_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n704_), .A2(new_n722_), .A3(new_n636_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n702_), .A2(new_n643_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n588_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT112), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n658_), .A2(new_n661_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n547_), .A2(new_n561_), .A3(new_n481_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n309_), .A2(new_n492_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n729_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n727_), .B2(new_n609_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n608_), .A2(new_n491_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n742_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n727_), .A2(new_n500_), .A3(new_n628_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n262_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n745_));
  INV_X1    g544(.A(G99gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT51), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n744_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n727_), .A2(new_n499_), .A3(new_n394_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n734_), .A2(new_n394_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G106gat), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT52), .B(new_n499_), .C1(new_n734_), .C2(new_n394_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n752_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NAND3_X1  g560(.A1(new_n429_), .A2(new_n588_), .A3(new_n628_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(KEYINPUT59), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n586_), .A2(new_n483_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n586_), .A2(new_n483_), .A3(new_n765_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n527_), .A2(new_n529_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n486_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n536_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n522_), .A4(new_n520_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n474_), .B1(new_n467_), .B2(new_n460_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n459_), .A2(new_n466_), .A3(new_n461_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n477_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n773_), .A2(new_n780_), .A3(new_n477_), .A4(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(KEYINPUT116), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT55), .B1(new_n530_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n770_), .A2(new_n486_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n536_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n536_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n782_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n782_), .B(KEYINPUT58), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n585_), .A3(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n481_), .A2(new_n774_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n789_), .A2(new_n798_), .A3(new_n536_), .A4(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n530_), .A2(new_n785_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n787_), .B1(new_n802_), .B2(new_n783_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n772_), .B1(new_n803_), .B2(new_n786_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n804_), .B2(new_n800_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n798_), .B1(new_n804_), .B2(KEYINPUT56), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n797_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n544_), .A2(new_n477_), .A3(new_n540_), .A4(new_n777_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n584_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n796_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n810_), .A2(KEYINPUT121), .B1(KEYINPUT57), .B2(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n796_), .B(new_n812_), .C1(new_n809_), .C2(KEYINPUT57), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n595_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n769_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT122), .B(new_n595_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n763_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(KEYINPUT120), .B2(new_n796_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n796_), .A2(KEYINPUT120), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(KEYINPUT57), .B2(new_n809_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n595_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n767_), .A2(new_n768_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n762_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n482_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G113gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n762_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n591_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1340gat));
  NAND3_X1  g631(.A1(new_n818_), .A2(new_n547_), .A3(new_n826_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  INV_X1    g633(.A(new_n762_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  AOI21_X1  g635(.A(G120gat), .B1(new_n547_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n836_), .B2(G120gat), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n835_), .B(new_n838_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT123), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(G1341gat));
  NAND3_X1  g640(.A1(new_n818_), .A2(new_n595_), .A3(new_n826_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G127gat), .ZN(new_n843_));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n829_), .A2(new_n844_), .A3(new_n595_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1342gat));
  NAND3_X1  g645(.A1(new_n818_), .A2(new_n585_), .A3(new_n826_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G134gat), .ZN(new_n848_));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n829_), .A2(new_n849_), .A3(new_n599_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n421_), .A2(new_n628_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n825_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n609_), .A2(new_n309_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G141gat), .B1(new_n856_), .B2(new_n481_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n854_), .A2(new_n264_), .A3(new_n591_), .A4(new_n855_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1344gat));
  OAI21_X1  g658(.A(G148gat), .B1(new_n856_), .B2(new_n546_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n854_), .A2(new_n265_), .A3(new_n547_), .A4(new_n855_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1345gat));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n856_), .B2(new_n561_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n854_), .A2(new_n595_), .A3(new_n855_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(new_n856_), .ZN(new_n868_));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n671_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n854_), .A2(new_n599_), .A3(new_n855_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n868_), .A2(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n608_), .A2(new_n588_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n628_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n636_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n591_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n810_), .A2(KEYINPUT121), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n813_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n561_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n824_), .B1(new_n882_), .B2(KEYINPUT122), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n814_), .A2(new_n815_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n878_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n873_), .B(new_n874_), .C1(new_n885_), .C2(new_n212_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n212_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n873_), .A2(new_n874_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n816_), .A2(new_n817_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(new_n888_), .C1(new_n889_), .C2(new_n878_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n885_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n886_), .A2(new_n890_), .A3(new_n891_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n547_), .A2(G176gat), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n825_), .A2(new_n394_), .A3(new_n876_), .A4(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n889_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n547_), .A3(new_n877_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n896_), .B2(new_n213_), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n329_), .A2(new_n331_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n595_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n877_), .B(new_n900_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n876_), .A2(new_n561_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n421_), .B(new_n902_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n206_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT125), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n901_), .A2(new_n904_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1350gat));
  OAI211_X1 g708(.A(new_n585_), .B(new_n877_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G190gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n895_), .A2(new_n877_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n599_), .A2(new_n332_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1351gat));
  AND2_X1   g713(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n852_), .B(new_n875_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n481_), .ZN(new_n919_));
  MUX2_X1   g718(.A(new_n917_), .B(new_n916_), .S(new_n919_), .Z(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n546_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(G204gat), .Z(G1353gat));
  OR2_X1    g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n918_), .A2(new_n561_), .ZN(new_n925_));
  MUX2_X1   g724(.A(new_n923_), .B(new_n924_), .S(new_n925_), .Z(G1354gat));
  INV_X1    g725(.A(new_n585_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT127), .B(G218gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n918_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n918_), .A2(new_n598_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(G1355gat));
endmodule


