//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n216_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(G92gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(G85gat), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n204_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(G92gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n216_), .A2(G85gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT9), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n208_), .A2(new_n209_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n223_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n211_), .A2(KEYINPUT8), .A3(new_n212_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n215_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G71gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G71gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G78gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G57gat), .A2(G64gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G57gat), .A2(G64gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT11), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n238_), .ZN(new_n244_));
  INV_X1    g043(.A(G78gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n235_), .A3(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(new_n241_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n242_), .B2(new_n238_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n233_), .A2(new_n235_), .A3(new_n245_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n231_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n215_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n247_), .A2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT66), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G120gat), .B(G148gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(G204gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT5), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT12), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(new_n231_), .B2(new_n252_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(KEYINPUT12), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n254_), .A2(new_n255_), .A3(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n269_), .A2(new_n271_), .A3(new_n258_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n257_), .A2(new_n259_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n261_), .B(new_n266_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n266_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n260_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT15), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G43gat), .B(G50gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(G29gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT68), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G29gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n298_), .A2(new_n294_), .A3(new_n287_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n286_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n296_), .A3(new_n288_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n287_), .B1(new_n298_), .B2(new_n294_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n254_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n297_), .A2(new_n299_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n231_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G232gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT34), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n305_), .B(new_n307_), .C1(KEYINPUT35), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT35), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT36), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G134gat), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n312_), .A2(new_n313_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n318_), .B(new_n314_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n321_), .A3(new_n313_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT37), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(KEYINPUT37), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n322_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n323_), .B(KEYINPUT37), .C1(new_n327_), .C2(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n255_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G15gat), .B(G22gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n333_));
  INV_X1    g132(.A(G8gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT71), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G8gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n333_), .A2(new_n335_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT14), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n339_), .B2(KEYINPUT14), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n332_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT73), .B(G1gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G8gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n332_), .B(new_n345_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n331_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G155gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G183gat), .B(G211gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT17), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n355_), .A2(KEYINPUT74), .A3(new_n356_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n350_), .A2(new_n358_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n329_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT76), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT76), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n285_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G85gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G134gat), .ZN(new_n374_));
  INV_X1    g173(.A(G127gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT80), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G127gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n374_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G113gat), .B(G120gat), .Z(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n378_), .A3(new_n374_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n381_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n382_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n379_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n394_), .B2(new_n390_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398_));
  INV_X1    g197(.A(G141gat), .ZN(new_n399_));
  INV_X1    g198(.A(G148gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G155gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n317_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n390_), .A3(new_n389_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n392_), .A2(KEYINPUT1), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n403_), .A2(new_n407_), .A3(new_n397_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT82), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n397_), .B(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n394_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n404_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n388_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n387_), .A2(new_n416_), .A3(new_n410_), .A4(new_n404_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT4), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n388_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n373_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n373_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G197gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT84), .B1(new_n432_), .B2(G204gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G211gat), .A2(G218gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G211gat), .A2(G218gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G211gat), .ZN(new_n439_));
  INV_X1    g238(.A(G218gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT85), .B1(new_n441_), .B2(new_n434_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT21), .B(new_n433_), .C1(new_n438_), .C2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G197gat), .B(G204gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n437_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(KEYINPUT85), .A3(new_n434_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n448_), .A2(KEYINPUT21), .ZN(new_n449_));
  INV_X1    g248(.A(new_n444_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(KEYINPUT21), .A3(new_n450_), .A4(new_n433_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n453_));
  AND2_X1   g252(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n454_));
  AND2_X1   g253(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n456_));
  OAI22_X1  g255(.A1(new_n453_), .A2(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT23), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT23), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G183gat), .A3(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  OR3_X1    g261(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n463_));
  INV_X1    g262(.A(G169gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n265_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT24), .A3(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .A4(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(G183gat), .A2(G190gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n471_));
  AND2_X1   g270(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n471_), .B(new_n265_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT22), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n464_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(G176gat), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n466_), .B1(new_n479_), .B2(new_n471_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n468_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n265_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT78), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(new_n470_), .A3(new_n466_), .A4(new_n474_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT79), .A3(new_n468_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n452_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n466_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n484_), .A2(KEYINPUT88), .A3(new_n466_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n470_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n468_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n494_), .A2(new_n449_), .A3(new_n451_), .A4(new_n445_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n495_), .A3(KEYINPUT20), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT19), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n483_), .A2(new_n487_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n445_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n498_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n452_), .A2(new_n468_), .A3(new_n493_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n503_), .A4(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT18), .B(G64gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G92gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT94), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(KEYINPUT94), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n503_), .B1(new_n517_), .B2(new_n504_), .ZN(new_n518_));
  AND4_X1   g317(.A1(KEYINPUT20), .A2(new_n488_), .A3(new_n495_), .A4(new_n503_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n514_), .B(new_n515_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n499_), .A2(new_n505_), .A3(KEYINPUT95), .A4(new_n509_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n512_), .A2(new_n520_), .A3(KEYINPUT27), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT27), .ZN(new_n523_));
  INV_X1    g322(.A(new_n510_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n509_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n404_), .A2(new_n410_), .A3(new_n529_), .A4(new_n416_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G22gat), .B(G50gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT28), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n532_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT87), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n452_), .B1(KEYINPUT29), .B2(new_n417_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G228gat), .A2(G233gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT86), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n417_), .A2(KEYINPUT29), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT83), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n417_), .A2(KEYINPUT83), .A3(KEYINPUT29), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n539_), .A3(new_n501_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n501_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT86), .ZN(new_n547_));
  INV_X1    g346(.A(new_n539_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n533_), .A2(KEYINPUT87), .A3(new_n534_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n540_), .A2(new_n545_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n537_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G71gat), .B(G99gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n486_), .A2(KEYINPUT79), .A3(new_n468_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT79), .B1(new_n486_), .B2(new_n468_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n560_), .A2(new_n561_), .A3(KEYINPUT30), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n387_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT30), .B1(new_n560_), .B2(new_n561_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n483_), .A2(new_n563_), .A3(new_n487_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n388_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G15gat), .B(G43gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT31), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n565_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n559_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n565_), .A2(new_n568_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n570_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n565_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n558_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n540_), .A2(new_n549_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n552_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n545_), .A4(new_n550_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n551_), .A2(new_n552_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n536_), .A3(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n555_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n555_), .B2(new_n584_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n431_), .B(new_n528_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n555_), .A2(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n590_));
  OR2_X1    g389(.A1(KEYINPUT90), .A2(KEYINPUT33), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n429_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n499_), .A2(new_n505_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n513_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT89), .A3(new_n510_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n420_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n418_), .A2(new_n422_), .A3(new_n419_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n372_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT91), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n597_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(KEYINPUT91), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n598_), .A2(new_n601_), .A3(new_n602_), .A4(new_n603_), .ZN(new_n604_));
  AND4_X1   g403(.A1(new_n590_), .A2(new_n592_), .A3(new_n595_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n509_), .A2(KEYINPUT32), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n499_), .A2(new_n505_), .A3(new_n606_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n425_), .A2(new_n426_), .A3(new_n373_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n608_), .B(new_n609_), .C1(new_n427_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n430_), .A2(KEYINPUT93), .A3(new_n609_), .A4(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n579_), .B(new_n588_), .C1(new_n605_), .C2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n587_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n347_), .A2(new_n306_), .A3(new_n348_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n306_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n342_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT14), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n345_), .B1(new_n625_), .B2(new_n332_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n348_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n304_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n347_), .A2(new_n306_), .A3(new_n348_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n618_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n464_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(new_n432_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n622_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n368_), .A2(new_n617_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n368_), .A2(new_n638_), .A3(KEYINPUT96), .A4(new_n617_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n333_), .A2(new_n338_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n430_), .B(KEYINPUT97), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n327_), .A2(new_n319_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n361_), .B(new_n652_), .C1(new_n587_), .C2(new_n616_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n622_), .A2(new_n630_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n633_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n622_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n285_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n431_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT99), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n647_), .A2(new_n649_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n650_), .A2(new_n661_), .A3(new_n662_), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n335_), .A2(new_n337_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n643_), .A2(new_n664_), .A3(new_n527_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G8gat), .B1(new_n659_), .B2(new_n528_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n667_));
  NOR2_X1   g466(.A1(KEYINPUT100), .A2(KEYINPUT39), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n665_), .A2(new_n669_), .A3(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n659_), .B2(new_n579_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT41), .Z(new_n676_));
  OR2_X1    g475(.A1(new_n639_), .A2(G15gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n579_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n659_), .B2(new_n588_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT101), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n639_), .A2(G22gat), .A3(new_n588_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(G1327gat));
  AOI21_X1  g484(.A(new_n651_), .B1(new_n587_), .B2(new_n616_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n361_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n285_), .A2(new_n637_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n430_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n617_), .B2(new_n329_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n329_), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT43), .B(new_n694_), .C1(new_n587_), .C2(new_n616_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n688_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT44), .Z(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n645_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n691_), .B1(new_n699_), .B2(G29gat), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n698_), .B2(new_n528_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n690_), .A2(new_n289_), .A3(new_n527_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT45), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n701_), .B(new_n703_), .C1(new_n705_), .C2(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(new_n579_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G43gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n689_), .A2(new_n579_), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n698_), .A2(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n698_), .B2(new_n588_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n588_), .A2(G50gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT103), .Z(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n689_), .B2(new_n717_), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n285_), .A2(new_n637_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n653_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n431_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n364_), .A2(new_n365_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n617_), .A3(new_n720_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n645_), .B1(new_n726_), .B2(KEYINPUT104), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(KEYINPUT104), .B2(new_n726_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n728_), .B2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n721_), .B2(new_n528_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT48), .Z(new_n731_));
  NOR3_X1   g530(.A1(new_n725_), .A2(G64gat), .A3(new_n528_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n721_), .B2(new_n579_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT49), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n232_), .A3(new_n710_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n721_), .B2(new_n588_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  INV_X1    g538(.A(new_n588_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n245_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n719_), .A2(new_n687_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n686_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT105), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n646_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT106), .Z(new_n747_));
  AND2_X1   g546(.A1(new_n696_), .A2(new_n743_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n431_), .A2(new_n224_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n745_), .B2(new_n527_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n219_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n218_), .A2(G92gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n528_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n748_), .B2(new_n754_), .ZN(G1337gat));
  NAND2_X1  g554(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n745_), .B(new_n710_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n696_), .A2(new_n710_), .A3(new_n743_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G99gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT107), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT107), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n756_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n762_), .B(new_n763_), .Z(G1338gat));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n740_), .B(new_n743_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G106gat), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n766_), .A2(new_n771_), .A3(new_n772_), .A4(G106gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n766_), .A2(new_n772_), .A3(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT109), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n767_), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n770_), .A2(new_n773_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n745_), .A2(new_n204_), .A3(new_n740_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n765_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n775_), .A2(new_n773_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT110), .B1(new_n767_), .B2(KEYINPUT52), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n769_), .B(new_n772_), .C1(new_n766_), .C2(G106gat), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n779_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT111), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(KEYINPUT53), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n782_), .A2(new_n790_), .ZN(G1339gat));
  NAND3_X1  g590(.A1(new_n646_), .A2(new_n586_), .A3(new_n528_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT118), .Z(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n618_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n633_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n628_), .A2(new_n619_), .A3(new_n629_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(KEYINPUT115), .A3(new_n633_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n656_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n282_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(KEYINPUT114), .B2(KEYINPUT56), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n254_), .A2(new_n255_), .A3(new_n272_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n272_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n258_), .B1(new_n807_), .B2(new_n269_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n274_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(new_n809_), .A3(new_n259_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n804_), .B1(new_n814_), .B2(new_n279_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816_));
  AND4_X1   g615(.A1(new_n258_), .A2(new_n269_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n811_), .A2(new_n259_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(KEYINPUT55), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(new_n279_), .C1(new_n819_), .C2(new_n812_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT114), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n815_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n280_), .A2(new_n279_), .A3(new_n260_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n637_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n657_), .A2(new_n278_), .A3(KEYINPUT112), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n803_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n794_), .B1(new_n829_), .B2(new_n652_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n827_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n820_), .B2(KEYINPUT114), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n815_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n651_), .C1(new_n833_), .C2(new_n803_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n266_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(KEYINPUT56), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n279_), .B1(new_n819_), .B2(new_n812_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT117), .A3(new_n822_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT56), .B(new_n279_), .C1(new_n819_), .C2(new_n812_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n838_), .A2(new_n840_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n802_), .A2(new_n825_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT58), .B1(new_n845_), .B2(new_n846_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n694_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n361_), .B1(new_n835_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n658_), .A2(new_n362_), .A3(new_n637_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT54), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n658_), .A2(new_n362_), .A3(new_n853_), .A4(new_n637_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n793_), .B1(new_n850_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n657_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n856_), .B(KEYINPUT59), .Z(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n637_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n858_), .B2(new_n658_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n658_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n856_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1341gat));
  NAND2_X1  g664(.A1(new_n687_), .A2(G127gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT119), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n856_), .A2(new_n687_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n858_), .A2(new_n868_), .B1(G127gat), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n856_), .B2(new_n652_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n858_), .A2(new_n694_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT121), .B(G134gat), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n850_), .A2(new_n855_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n877_), .A2(new_n585_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n878_), .A2(new_n528_), .A3(new_n646_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n657_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n285_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n687_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n879_), .B2(new_n652_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n694_), .A2(new_n317_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n879_), .B2(new_n888_), .ZN(G1347gat));
  AND2_X1   g688(.A1(new_n586_), .A2(new_n527_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n877_), .A2(new_n657_), .A3(new_n645_), .A4(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT122), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n646_), .B1(new_n850_), .B2(new_n855_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n657_), .A4(new_n890_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(G169gat), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n892_), .A2(new_n895_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .A4(G169gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT123), .B1(new_n896_), .B2(KEYINPUT62), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n896_), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n899_), .A2(new_n903_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n893_), .A2(new_n890_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n908_), .B(new_n657_), .C1(new_n473_), .C2(new_n472_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(G1348gat));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n658_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n265_), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n687_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  INV_X1    g714(.A(G183gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n913_), .B2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n914_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(KEYINPUT125), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n907_), .B2(new_n694_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n652_), .B1(new_n456_), .B2(new_n455_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n907_), .B2(new_n921_), .ZN(G1351gat));
  NOR2_X1   g721(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT126), .B(G197gat), .Z(new_n924_));
  AND4_X1   g723(.A1(new_n431_), .A2(new_n877_), .A3(new_n585_), .A4(new_n527_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n657_), .ZN(new_n926_));
  MUX2_X1   g725(.A(new_n923_), .B(new_n924_), .S(new_n926_), .Z(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n285_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n439_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n925_), .A2(new_n687_), .A3(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n439_), .ZN(new_n933_));
  OR3_X1    g732(.A1(new_n932_), .A2(KEYINPUT127), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n925_), .A2(new_n687_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n935_), .A2(new_n930_), .A3(new_n439_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n932_), .B2(new_n933_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n934_), .A2(new_n936_), .A3(new_n937_), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n925_), .B2(new_n652_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n925_), .A2(new_n329_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(G218gat), .B2(new_n940_), .ZN(G1355gat));
endmodule


