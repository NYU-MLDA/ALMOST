//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT83), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT22), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(G169gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT80), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214_));
  AOI21_X1  g013(.A(G176gat), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n212_), .A2(new_n215_), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT81), .B1(new_n217_), .B2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n224_), .A2(new_n221_), .A3(G183gat), .A4(G190gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n219_), .A2(new_n220_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n216_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n234_), .B2(KEYINPUT78), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(G190gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(KEYINPUT26), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(KEYINPUT26), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n238_), .B1(new_n242_), .B2(new_n236_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n208_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(KEYINPUT24), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n222_), .ZN(new_n250_));
  OR3_X1    g049(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n244_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n228_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n207_), .B1(new_n255_), .B2(KEYINPUT84), .ZN(new_n256_));
  AND2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n224_), .B1(new_n257_), .B2(new_n221_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n217_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n217_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n258_), .A2(new_n259_), .B1(new_n260_), .B2(new_n218_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n227_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n263_), .A2(new_n216_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT30), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n207_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G113gat), .B(G120gat), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G113gat), .B(G120gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(KEYINPUT85), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n275_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT31), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n270_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n268_), .A2(new_n281_), .A3(new_n269_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G155gat), .B(G162gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n288_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G141gat), .B(G148gat), .Z(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n296_), .B(new_n297_), .C1(KEYINPUT1), .C2(new_n287_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G197gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(KEYINPUT21), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT87), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n312_), .A2(new_n307_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n304_), .A2(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n303_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n325_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n302_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(new_n302_), .A3(new_n327_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n332_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n328_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n286_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n280_), .A2(new_n299_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT95), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n280_), .A2(new_n299_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n274_), .A2(new_n276_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n277_), .A2(new_n279_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n341_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT0), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G57gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n361_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n362_), .A2(G85gat), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(G85gat), .B1(new_n362_), .B2(new_n363_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n355_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n371_));
  AND2_X1   g170(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n372_));
  OAI22_X1  g171(.A1(new_n371_), .A2(new_n366_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT97), .ZN(new_n375_));
  INV_X1    g174(.A(new_n346_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n348_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n344_), .A2(KEYINPUT97), .A3(new_n346_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n353_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n366_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT98), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT98), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n366_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n351_), .A2(new_n353_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT99), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n381_), .A2(new_n384_), .A3(new_n387_), .A4(new_n383_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n374_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n310_), .A2(new_n315_), .B1(new_n318_), .B2(new_n317_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT89), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT89), .B1(new_n239_), .B2(new_n241_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n234_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n248_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n242_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT89), .ZN(new_n401_));
  INV_X1    g200(.A(new_n234_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT90), .A3(new_n248_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n261_), .A2(new_n251_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n398_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n245_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n247_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n410_), .A2(new_n411_), .B1(new_n262_), .B2(new_n250_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(KEYINPUT91), .A3(new_n247_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n392_), .B1(new_n407_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n320_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n391_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT92), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT94), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n421_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n391_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n264_), .B2(new_n392_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n403_), .A2(new_n248_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n405_), .B1(new_n429_), .B2(new_n393_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n430_), .A2(new_n404_), .B1(new_n413_), .B2(new_n412_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n431_), .B2(new_n392_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n391_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n418_), .A2(new_n425_), .A3(new_n427_), .A4(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n417_), .A2(KEYINPUT92), .B1(new_n432_), .B2(new_n433_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n425_), .B1(new_n437_), .B2(new_n427_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n357_), .A2(new_n367_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n371_), .A2(new_n366_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT32), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n424_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n264_), .B2(new_n392_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n433_), .B(new_n447_), .C1(new_n431_), .C2(new_n392_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n407_), .A2(new_n392_), .A3(new_n414_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n254_), .B2(new_n320_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n433_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT101), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT101), .B(new_n433_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n445_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n445_), .B(KEYINPUT100), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n437_), .A2(new_n427_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n443_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n389_), .A2(new_n439_), .B1(new_n440_), .B2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n440_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n340_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n418_), .A2(new_n427_), .A3(new_n434_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n424_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT27), .B1(new_n463_), .B2(new_n435_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n424_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n465_), .A2(KEYINPUT27), .A3(new_n435_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT103), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT27), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT103), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(KEYINPUT27), .A3(new_n435_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n338_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n339_), .A2(new_n285_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n443_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n461_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT10), .B(G99gat), .Z(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G85gat), .B(G92gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT9), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT6), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n484_), .A2(new_n486_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  OR3_X1    g292(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n485_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n495_), .B2(new_n485_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n492_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT65), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(new_n492_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G43gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G43gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n504_), .B(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT71), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n503_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(KEYINPUT71), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n506_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(G50gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n511_), .A2(KEYINPUT15), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT15), .B1(new_n511_), .B2(new_n514_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n500_), .B(new_n502_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT69), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT34), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n511_), .A2(new_n514_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(new_n523_), .B2(new_n499_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT70), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n527_), .A3(KEYINPUT73), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT72), .B(new_n522_), .C1(new_n523_), .C2(new_n499_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n524_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n518_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n530_), .A2(new_n531_), .B1(new_n526_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT36), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n481_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n535_), .A2(new_n526_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n531_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT73), .B1(new_n518_), .B2(new_n527_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(KEYINPUT74), .A3(new_n540_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n530_), .A2(new_n531_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n541_), .B1(new_n552_), .B2(new_n545_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n550_), .A2(new_n551_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G1gat), .ZN(new_n557_));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT14), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT75), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n560_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G1gat), .B(G8gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G71gat), .B(G78gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(KEYINPUT11), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n568_), .B(new_n573_), .Z(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n229_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G211gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n566_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n523_), .A2(new_n584_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT76), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT76), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n585_), .A2(new_n591_), .A3(new_n586_), .A4(new_n588_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n523_), .B(new_n584_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n586_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G169gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n306_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT77), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n590_), .A2(new_n603_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n499_), .A2(new_n573_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT12), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n499_), .A2(new_n573_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT64), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n500_), .A2(KEYINPUT12), .A3(new_n502_), .A4(new_n573_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n608_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n615_), .B2(new_n606_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT67), .ZN(new_n619_));
  XOR2_X1   g418(.A(G120gat), .B(G148gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n623_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(new_n616_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT13), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(KEYINPUT13), .A3(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT68), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(KEYINPUT68), .A3(new_n630_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n605_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n556_), .A2(new_n583_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n480_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n443_), .B(KEYINPUT104), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n557_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  INV_X1    g439(.A(new_n550_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n479_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n631_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n605_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n583_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n478_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n640_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT105), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n467_), .A2(new_n472_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n480_), .A2(new_n636_), .A3(new_n558_), .A4(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n652_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G8gat), .B1(new_n648_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT39), .B(G8gat), .C1(new_n648_), .C2(new_n656_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT107), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n655_), .A2(new_n659_), .A3(new_n663_), .A4(new_n660_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n662_), .A2(KEYINPUT40), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT40), .B1(new_n662_), .B2(new_n664_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n648_), .B2(new_n286_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  INV_X1    g468(.A(new_n637_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n286_), .A2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n670_), .B2(new_n671_), .ZN(G1326gat));
  OAI21_X1  g471(.A(G22gat), .B1(new_n648_), .B2(new_n339_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n339_), .A2(G22gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n670_), .B2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n479_), .A2(new_n550_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n645_), .A2(new_n583_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n443_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n477_), .A2(new_n478_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n461_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n556_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n550_), .A2(new_n551_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n554_), .A2(new_n555_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n443_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n461_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT43), .B1(new_n692_), .B2(KEYINPUT109), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n687_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n682_), .B(KEYINPUT43), .C1(new_n685_), .C2(new_n686_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(KEYINPUT44), .A3(new_n678_), .A4(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(G29gat), .A3(new_n638_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n685_), .B2(new_n682_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT109), .B1(new_n692_), .B2(KEYINPUT108), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n695_), .B(new_n678_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n681_), .B1(new_n697_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n696_), .A2(new_n652_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n703_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n679_), .A2(G36gat), .A3(new_n656_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n703_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n696_), .A2(new_n652_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G36gat), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(KEYINPUT46), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1329gat));
  XOR2_X1   g516(.A(KEYINPUT110), .B(G43gat), .Z(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n679_), .B2(new_n286_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n696_), .A2(G43gat), .A3(new_n285_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n712_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n680_), .B2(new_n338_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n696_), .A2(G50gat), .A3(new_n338_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n703_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n643_), .A2(new_n644_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n690_), .A2(new_n727_), .A3(new_n646_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n480_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n638_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT111), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n633_), .A2(new_n634_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n605_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n646_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n642_), .A2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n361_), .A3(new_n478_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n731_), .A2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n735_), .B2(new_n656_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  INV_X1    g538(.A(new_n729_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n656_), .A2(G64gat), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT112), .Z(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n740_), .B2(new_n742_), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n744_), .A3(new_n285_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n735_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n285_), .ZN(new_n747_));
  XOR2_X1   g546(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n747_), .A2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT114), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n735_), .B2(new_n339_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n339_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n740_), .B2(new_n757_), .ZN(G1335gat));
  OAI21_X1  g557(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n694_), .A2(KEYINPUT116), .A3(new_n695_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n727_), .A2(new_n583_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n487_), .B1(new_n764_), .B2(new_n443_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n733_), .A2(new_n583_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n677_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n638_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n767_), .A2(G85gat), .A3(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n765_), .A2(new_n769_), .ZN(G1336gat));
  OAI21_X1  g569(.A(new_n488_), .B1(new_n767_), .B2(new_n656_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT117), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n656_), .A2(new_n488_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n764_), .B2(new_n773_), .ZN(G1337gat));
  NAND4_X1  g573(.A1(new_n761_), .A2(new_n285_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G99gat), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n677_), .A2(new_n766_), .A3(new_n285_), .A4(new_n482_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT51), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1338gat));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n483_), .B1(new_n783_), .B2(KEYINPUT52), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n763_), .A2(new_n338_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n759_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT119), .A3(new_n787_), .ZN(new_n788_));
  OAI221_X1 g587(.A(new_n784_), .B1(new_n783_), .B2(KEYINPUT52), .C1(new_n759_), .C2(new_n785_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n767_), .A2(G106gat), .A3(new_n339_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT118), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n788_), .A2(new_n791_), .A3(new_n794_), .A4(new_n789_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  XNOR2_X1  g595(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n652_), .A2(new_n768_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT15), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n523_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n566_), .B1(new_n802_), .B2(new_n515_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n803_), .B2(new_n587_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n585_), .A2(KEYINPUT121), .A3(new_n588_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n586_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n593_), .A2(new_n594_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n600_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n590_), .A2(new_n599_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n612_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n614_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n609_), .A2(KEYINPUT55), .A3(new_n612_), .A4(new_n613_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n625_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n626_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n810_), .A2(new_n818_), .A3(KEYINPUT58), .A4(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  INV_X1    g622(.A(new_n821_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n808_), .B(new_n809_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n553_), .A2(KEYINPUT74), .B1(new_n536_), .B2(new_n543_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT37), .B1(new_n827_), .B2(new_n542_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n689_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n822_), .B(new_n826_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n808_), .A2(new_n627_), .A3(new_n809_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n602_), .A2(new_n626_), .A3(new_n604_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n815_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n835_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n625_), .B(new_n837_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n832_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n831_), .B1(new_n840_), .B2(new_n641_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n833_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT57), .B(new_n550_), .C1(new_n842_), .C2(new_n832_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n830_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n646_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n644_), .A2(new_n631_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n556_), .A2(new_n583_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n556_), .A2(new_n849_), .A3(new_n583_), .A4(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n799_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n797_), .B1(new_n852_), .B2(new_n473_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n844_), .A2(new_n646_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n473_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n799_), .A4(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT124), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n857_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n852_), .A2(new_n473_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n854_), .A2(new_n855_), .A3(new_n799_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n861_), .B(new_n862_), .C1(new_n863_), .C2(new_n797_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n864_), .A3(new_n644_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G113gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n863_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n867_), .A2(G113gat), .A3(new_n605_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1340gat));
  NOR2_X1   g668(.A1(new_n643_), .A2(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n863_), .B1(KEYINPUT60), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n732_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n861_), .B1(new_n863_), .B2(new_n797_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G120gat), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(G1341gat));
  AOI21_X1  g674(.A(G127gat), .B1(new_n863_), .B2(new_n583_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n859_), .A2(new_n864_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n583_), .A2(G127gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT125), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1342gat));
  NAND3_X1  g679(.A1(new_n859_), .A2(new_n864_), .A3(new_n690_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G134gat), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n867_), .A2(G134gat), .A3(new_n550_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  INV_X1    g683(.A(new_n475_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n854_), .A2(new_n885_), .A3(new_n799_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n644_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n732_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n583_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n886_), .B2(new_n641_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n690_), .A2(G162gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT126), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n886_), .B2(new_n896_), .ZN(G1347gat));
  NAND3_X1  g696(.A1(new_n652_), .A2(new_n473_), .A3(new_n768_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n854_), .A2(new_n605_), .A3(new_n898_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n899_), .A2(new_n208_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n408_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n901_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n854_), .A2(new_n898_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906_), .B2(new_n631_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n732_), .A2(G176gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n583_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n402_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n229_), .B2(new_n910_), .ZN(G1350gat));
  NAND4_X1  g711(.A1(new_n906_), .A2(new_n400_), .A3(new_n401_), .A4(new_n641_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n854_), .A2(new_n556_), .A3(new_n898_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n237_), .ZN(G1351gat));
  NOR4_X1   g714(.A1(new_n854_), .A2(new_n443_), .A3(new_n885_), .A4(new_n656_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n644_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT127), .B(G197gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n732_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n583_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n916_), .A2(new_n927_), .A3(new_n641_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n916_), .A2(new_n690_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n927_), .ZN(G1355gat));
endmodule


