//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT23), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n202_), .B(new_n205_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n204_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n211_), .A2(KEYINPUT83), .A3(KEYINPUT26), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT83), .B1(new_n211_), .B2(KEYINPUT26), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n222_), .B(new_n223_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n212_), .A2(new_n207_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT86), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT31), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G15gat), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT85), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n230_), .B2(KEYINPUT86), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  INV_X1    g044(.A(G120gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT87), .B(G113gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n244_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n237_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n235_), .A2(new_n236_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT90), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT2), .Z(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n257_), .B(new_n258_), .C1(new_n260_), .C2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n261_), .B(KEYINPUT89), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n258_), .B(KEYINPUT1), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n259_), .B1(new_n256_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n249_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT102), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n249_), .B(new_n268_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n270_), .B(new_n273_), .C1(new_n274_), .C2(new_n269_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n271_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G85gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G57gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n275_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n268_), .A2(KEYINPUT29), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT28), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G22gat), .B(G50gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n268_), .A2(KEYINPUT29), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292_));
  INV_X1    g091(.A(G197gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(G204gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(G197gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT21), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT93), .B1(new_n295_), .B2(G197gat), .ZN(new_n298_));
  MUX2_X1   g097(.A(new_n298_), .B(KEYINPUT93), .S(new_n294_), .Z(new_n299_));
  OAI211_X1 g098(.A(new_n292_), .B(new_n297_), .C1(new_n299_), .C2(KEYINPUT21), .ZN(new_n300_));
  INV_X1    g099(.A(new_n292_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(KEYINPUT21), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n291_), .A2(KEYINPUT92), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT91), .B(G228gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G78gat), .B(G106gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n304_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n290_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n254_), .A2(new_n286_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT98), .ZN(new_n313_));
  INV_X1    g112(.A(new_n202_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n203_), .B(KEYINPUT96), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n204_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n214_), .B1(new_n212_), .B2(new_n207_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT97), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n216_), .B(KEYINPUT95), .Z(new_n319_));
  AOI21_X1  g118(.A(new_n220_), .B1(new_n319_), .B2(new_n219_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G190gat), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n209_), .A2(new_n212_), .B1(new_n222_), .B2(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n316_), .A2(new_n318_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n303_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n313_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n316_), .A2(new_n318_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n320_), .A2(new_n322_), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT98), .B(new_n303_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n228_), .A3(new_n215_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n325_), .A2(new_n328_), .A3(KEYINPUT20), .A4(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT99), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n229_), .A2(new_n303_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n323_), .A2(new_n324_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT20), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n333_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT99), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n341_), .A3(new_n334_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT101), .ZN(new_n345_));
  XOR2_X1   g144(.A(G64gat), .B(G92gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n336_), .A2(new_n340_), .A3(new_n349_), .A4(new_n342_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT27), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n339_), .A2(new_n333_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n334_), .B2(new_n330_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n350_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n356_), .A2(new_n352_), .A3(KEYINPUT27), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n312_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n285_), .B(KEYINPUT33), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n270_), .B1(new_n274_), .B2(new_n269_), .ZN(new_n361_));
  OAI221_X1 g160(.A(new_n283_), .B1(new_n274_), .B2(new_n272_), .C1(new_n361_), .C2(new_n276_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n360_), .A2(new_n351_), .A3(new_n362_), .A4(new_n352_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n355_), .A2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n366_), .B(new_n286_), .C1(new_n365_), .C2(new_n343_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT103), .B1(new_n368_), .B2(new_n310_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT103), .ZN(new_n370_));
  AOI211_X1 g169(.A(new_n370_), .B(new_n311_), .C1(new_n363_), .C2(new_n367_), .ZN(new_n371_));
  NOR4_X1   g170(.A1(new_n353_), .A2(new_n357_), .A3(new_n286_), .A4(new_n310_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n254_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n359_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT7), .ZN(new_n378_));
  INV_X1    g177(.A(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(G106gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G99gat), .A2(G106gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n381_), .A2(new_n384_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G85gat), .A2(G92gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G85gat), .A2(G92gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT8), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(KEYINPUT8), .A3(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(KEYINPUT10), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G99gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(G106gat), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(new_n385_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT9), .B1(new_n388_), .B2(new_n389_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT66), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G85gat), .A2(G92gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT9), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n404_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT67), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n399_), .A2(new_n400_), .A3(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n407_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n395_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(G57gat), .A2(G64gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G57gat), .A2(G64gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT11), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G78gat), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT11), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n422_), .A3(new_n417_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n377_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n427_));
  NAND2_X1  g226(.A1(G230gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n387_), .A2(KEYINPUT8), .A3(new_n390_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT8), .B1(new_n387_), .B2(new_n390_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND4_X1   g232(.A1(new_n413_), .A2(new_n401_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n413_), .B1(new_n412_), .B2(new_n407_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n425_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT69), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n426_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT70), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n426_), .A2(new_n430_), .A3(new_n443_), .A4(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n425_), .B(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT68), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n411_), .A2(new_n414_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n425_), .A4(new_n433_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n425_), .B1(new_n448_), .B2(new_n433_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n429_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT5), .B(G176gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(new_n295_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G120gat), .B(G148gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n458_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n461_));
  OR3_X1    g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT71), .ZN(new_n463_));
  OAI22_X1  g262(.A1(new_n459_), .A2(new_n460_), .B1(new_n463_), .B2(KEYINPUT13), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT77), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G1gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n473_), .A3(G8gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT14), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n474_), .B2(KEYINPUT14), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n469_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n469_), .B(new_n479_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n468_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT79), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n489_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n467_), .B(KEYINPUT80), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n486_), .B(KEYINPUT15), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n493_), .B(new_n494_), .C1(new_n483_), .C2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT79), .B(new_n468_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n492_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT81), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(KEYINPUT81), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n499_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n492_), .A2(new_n497_), .A3(new_n498_), .A4(new_n503_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT82), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n506_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n466_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n415_), .A2(new_n486_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n436_), .A2(new_n495_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n518_), .A2(KEYINPUT35), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT74), .B1(new_n518_), .B2(KEYINPUT35), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n515_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT75), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT75), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n515_), .A2(new_n516_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n519_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n525_), .B2(new_n519_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n523_), .B(new_n524_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(KEYINPUT36), .A3(new_n534_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT76), .A3(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(KEYINPUT76), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(KEYINPUT76), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n483_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n425_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G211gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT16), .B(G183gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n549_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n555_), .B2(new_n549_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n546_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n375_), .A2(new_n514_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT104), .ZN(new_n562_));
  INV_X1    g361(.A(new_n471_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n473_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n562_), .B(new_n286_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT38), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n375_), .A2(new_n540_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT105), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n569_), .A2(new_n558_), .A3(new_n514_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(new_n286_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n470_), .B2(new_n571_), .ZN(G1324gat));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n358_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n562_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n569_), .A2(new_n558_), .A3(new_n514_), .A4(new_n574_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(G8gat), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n576_), .B2(G8gat), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n575_), .B(new_n581_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(G1325gat));
  INV_X1    g384(.A(G15gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n562_), .A2(new_n586_), .A3(new_n374_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n570_), .A2(new_n374_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n588_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT41), .B1(new_n588_), .B2(G15gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n589_), .B2(new_n590_), .ZN(G1326gat));
  NOR2_X1   g390(.A1(new_n310_), .A2(G22gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT107), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n562_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n570_), .A2(new_n311_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT42), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n595_), .A2(new_n596_), .A3(G22gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n595_), .B2(G22gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(G1327gat));
  NOR2_X1   g398(.A1(new_n540_), .A2(new_n558_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n375_), .A2(new_n514_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n286_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n368_), .A2(new_n310_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n370_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n368_), .A2(KEYINPUT103), .A3(new_n310_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n286_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n358_), .A2(new_n606_), .A3(new_n311_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n608_), .A2(new_n254_), .B1(new_n358_), .B2(new_n312_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n546_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT43), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT43), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n375_), .A2(new_n612_), .A3(new_n546_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n514_), .A2(new_n559_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT108), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(KEYINPUT44), .A3(new_n616_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n620_), .A2(new_n606_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n602_), .B1(new_n623_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g423(.A(KEYINPUT111), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT110), .B1(new_n625_), .B2(KEYINPUT46), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n574_), .A3(new_n621_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G36gat), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT109), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n601_), .A2(new_n629_), .A3(new_n630_), .A4(new_n574_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n375_), .A2(new_n630_), .A3(new_n514_), .A4(new_n600_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT109), .B1(new_n632_), .B2(new_n358_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n631_), .A2(KEYINPUT45), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT45), .B1(new_n631_), .B2(new_n633_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n626_), .B1(new_n628_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT110), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n628_), .A2(new_n638_), .A3(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n625_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n619_), .A2(G43gat), .A3(new_n374_), .A4(new_n621_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n601_), .A2(new_n374_), .ZN(new_n644_));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT112), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n644_), .A2(KEYINPUT112), .A3(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g448(.A(G50gat), .B1(new_n601_), .B2(new_n311_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n620_), .A2(new_n310_), .A3(new_n622_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g451(.A1(new_n465_), .A2(new_n512_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n609_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n560_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT113), .ZN(new_n657_));
  AOI21_X1  g456(.A(G57gat), .B1(new_n657_), .B2(new_n286_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n654_), .A2(new_n559_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n569_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(new_n286_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n658_), .B1(new_n661_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g461(.A(G64gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n660_), .B2(new_n574_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT48), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n663_), .A3(new_n574_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1333gat));
  INV_X1    g467(.A(G71gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n660_), .B2(new_n374_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT49), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n657_), .A2(new_n669_), .A3(new_n374_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1334gat));
  INV_X1    g473(.A(G78gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n660_), .B2(new_n311_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT50), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n657_), .A2(new_n675_), .A3(new_n311_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1335gat));
  AND2_X1   g479(.A1(new_n655_), .A2(new_n600_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G85gat), .B1(new_n681_), .B2(new_n286_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n558_), .B(new_n654_), .C1(new_n611_), .C2(new_n613_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n286_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n684_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g484(.A(G92gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n683_), .B2(new_n574_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n681_), .A2(new_n574_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT114), .Z(G1337gat));
  AOI21_X1  g489(.A(new_n379_), .B1(new_n683_), .B2(new_n374_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n254_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n681_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g493(.A1(new_n681_), .A2(new_n380_), .A3(new_n311_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n683_), .A2(new_n311_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G106gat), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT52), .B(new_n380_), .C1(new_n683_), .C2(new_n311_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT53), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT53), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n695_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1339gat));
  NOR2_X1   g503(.A1(new_n574_), .A2(new_n606_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n254_), .A2(new_n311_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT55), .B1(new_n442_), .B2(new_n444_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n440_), .B1(new_n452_), .B2(new_n376_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n429_), .B1(new_n451_), .B2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n426_), .A2(new_n430_), .A3(KEYINPUT55), .A4(new_n440_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n458_), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT56), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT116), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT56), .B(new_n458_), .C1(new_n708_), .C2(new_n712_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n460_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n708_), .A2(new_n712_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n458_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n512_), .A4(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT117), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n493_), .B1(new_n483_), .B2(new_n496_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n494_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n487_), .A2(new_n489_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n503_), .B(new_n725_), .C1(new_n494_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n511_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n509_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT116), .B1(new_n713_), .B2(new_n714_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n460_), .B1(new_n731_), .B2(new_n717_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n512_), .A4(new_n721_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n730_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n540_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n715_), .A2(new_n717_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n719_), .A3(new_n729_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT118), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT58), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT58), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n741_), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n546_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n540_), .A3(KEYINPUT57), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n743_), .A2(new_n546_), .A3(KEYINPUT119), .A4(new_n745_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n738_), .A2(new_n748_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n559_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n542_), .A2(new_n465_), .A3(new_n558_), .A4(new_n545_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n753_), .A2(new_n512_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n753_), .B2(new_n512_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n707_), .B1(new_n752_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G113gat), .B1(new_n759_), .B2(new_n512_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n751_), .A2(new_n559_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT59), .B1(new_n761_), .B2(new_n707_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n749_), .A2(new_n746_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(new_n735_), .B2(new_n540_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n559_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n758_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT59), .ZN(new_n767_));
  INV_X1    g566(.A(new_n707_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(new_n513_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n760_), .B1(new_n771_), .B2(G113gat), .ZN(G1340gat));
  OAI211_X1 g571(.A(new_n466_), .B(new_n769_), .C1(new_n759_), .C2(new_n767_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT120), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n762_), .A2(new_n775_), .A3(new_n466_), .A4(new_n769_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(G120gat), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n246_), .B1(new_n465_), .B2(KEYINPUT60), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n759_), .B(new_n778_), .C1(KEYINPUT60), .C2(new_n246_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(KEYINPUT121), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1341gat));
  NAND4_X1  g583(.A1(new_n762_), .A2(G127gat), .A3(new_n558_), .A4(new_n769_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n759_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n559_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(G127gat), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT122), .Z(G1342gat));
  AOI21_X1  g588(.A(G134gat), .B1(new_n759_), .B2(new_n539_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n770_), .A2(new_n610_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g591(.A1(new_n761_), .A2(new_n374_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n311_), .A3(new_n705_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n513_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT123), .B(G141gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1344gat));
  NOR2_X1   g596(.A1(new_n794_), .A2(new_n465_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT124), .B(G148gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1345gat));
  NOR2_X1   g599(.A1(new_n794_), .A2(new_n559_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT61), .B(G155gat), .Z(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1346gat));
  NOR2_X1   g602(.A1(new_n794_), .A2(new_n540_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(G162gat), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n794_), .A2(new_n610_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(G162gat), .B2(new_n806_), .ZN(G1347gat));
  NOR2_X1   g606(.A1(new_n358_), .A2(new_n286_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n766_), .A2(new_n706_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n512_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G169gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT62), .ZN(new_n813_));
  INV_X1    g612(.A(new_n315_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n811_), .ZN(G1348gat));
  AOI21_X1  g614(.A(G176gat), .B1(new_n810_), .B2(new_n466_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n374_), .A2(new_n808_), .ZN(new_n817_));
  NOR4_X1   g616(.A1(new_n761_), .A2(new_n204_), .A3(new_n311_), .A4(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n466_), .B2(new_n818_), .ZN(G1349gat));
  NOR3_X1   g618(.A1(new_n809_), .A2(new_n559_), .A3(new_n222_), .ZN(new_n820_));
  OR4_X1    g619(.A1(new_n559_), .A2(new_n761_), .A3(new_n311_), .A4(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n210_), .ZN(G1350gat));
  OAI21_X1  g621(.A(G190gat), .B1(new_n809_), .B2(new_n610_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n539_), .A2(new_n321_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n809_), .B2(new_n824_), .ZN(G1351gat));
  NAND3_X1  g624(.A1(new_n793_), .A2(new_n311_), .A3(new_n808_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT125), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n793_), .A2(new_n828_), .A3(new_n311_), .A4(new_n808_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT126), .B(G197gat), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n512_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n830_), .B2(new_n512_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1352gat));
  AOI21_X1  g633(.A(new_n465_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT127), .B(G204gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1353gat));
  XNOR2_X1  g636(.A(KEYINPUT63), .B(G211gat), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n559_), .B(new_n838_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n558_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(G1354gat));
  AOI21_X1  g641(.A(G218gat), .B1(new_n830_), .B2(new_n539_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n610_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(G218gat), .B2(new_n844_), .ZN(G1355gat));
endmodule


