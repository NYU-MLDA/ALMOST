//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n212_), .A2(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT82), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n209_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT92), .B1(new_n209_), .B2(KEYINPUT24), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G183gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n229_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n212_), .A2(new_n214_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n218_), .B1(new_n226_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(G197gat), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(G197gat), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .A4(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n240_), .A2(G197gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(G204gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT21), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G218gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G211gat), .ZN(new_n251_));
  INV_X1    g050(.A(G211gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G218gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT88), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT88), .B1(new_n251_), .B2(new_n253_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n246_), .B(new_n249_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n253_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n241_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT88), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT21), .A4(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n202_), .B1(new_n238_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT22), .B1(new_n268_), .B2(new_n205_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n269_), .B(new_n207_), .C1(new_n268_), .C2(new_n204_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n216_), .A2(KEYINPUT81), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT81), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n211_), .B(new_n213_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n270_), .B(new_n209_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n222_), .A2(new_n234_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT24), .A4(new_n209_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n231_), .B1(new_n274_), .B2(KEYINPUT26), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n228_), .A2(KEYINPUT80), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n227_), .A3(G183gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n284_), .A3(new_n229_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n277_), .B1(new_n280_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n256_), .A2(new_n262_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n264_), .A2(new_n267_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n278_), .B(new_n279_), .C1(new_n281_), .C2(new_n285_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n263_), .A2(new_n293_), .A3(new_n277_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n225_), .A2(new_n236_), .B1(new_n217_), .B2(new_n210_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n202_), .B1(new_n295_), .B2(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n267_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n264_), .A2(KEYINPUT93), .A3(new_n289_), .A4(new_n267_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G8gat), .B(G36gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n292_), .A2(new_n299_), .A3(new_n300_), .A4(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n294_), .A2(new_n296_), .A3(new_n267_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n267_), .B1(new_n264_), .B2(new_n289_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(KEYINPUT98), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n306_), .A2(KEYINPUT98), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT27), .B(new_n305_), .C1(new_n310_), .C2(new_n304_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n299_), .A2(new_n300_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n288_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n293_), .A2(new_n277_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT93), .B1(new_n316_), .B2(new_n267_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n305_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n311_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G155gat), .ZN(new_n324_));
  INV_X1    g123(.A(G162gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT85), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT85), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(G155gat), .B2(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(G141gat), .ZN(new_n333_));
  INV_X1    g132(.A(G148gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT3), .ZN(new_n335_));
  AND3_X1   g134(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n332_), .A2(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n339_), .A2(KEYINPUT86), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n330_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n334_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n340_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n326_), .A2(new_n328_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G155gat), .A3(G162gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n345_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT29), .B1(new_n343_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n352_), .A2(new_n288_), .B1(KEYINPUT89), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT90), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n356_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G22gat), .B(G50gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n343_), .A2(new_n351_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT28), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n366_), .A3(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n353_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n360_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n357_), .A2(new_n358_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n361_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n361_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n323_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT84), .B(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n287_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G127gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(G134gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(G134gat), .ZN(new_n385_));
  INV_X1    g184(.A(G113gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(G120gat), .ZN(new_n387_));
  INV_X1    g186(.A(G120gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(G113gat), .ZN(new_n389_));
  OAI22_X1  g188(.A1(new_n384_), .A2(new_n385_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n382_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT30), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n395_), .A2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n390_), .A2(new_n393_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n335_), .A2(new_n332_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n336_), .A2(new_n337_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n342_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n330_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n326_), .A2(new_n347_), .A3(new_n328_), .A4(new_n349_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n406_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n405_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n394_), .B1(new_n343_), .B2(new_n351_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n411_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT4), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n405_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G85gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT0), .B(G57gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n421_), .A2(new_n426_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n422_), .A2(new_n427_), .B1(new_n420_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n378_), .A2(new_n404_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n377_), .A2(new_n429_), .A3(new_n321_), .A4(new_n311_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n318_), .A2(new_n305_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n428_), .A2(new_n435_), .A3(new_n420_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n428_), .B2(new_n420_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT97), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n420_), .A2(KEYINPUT33), .A3(new_n421_), .A4(new_n426_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n428_), .A2(KEYINPUT94), .A3(KEYINPUT33), .A4(new_n420_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n419_), .B(new_n405_), .C1(KEYINPUT4), .C2(new_n417_), .ZN(new_n444_));
  AND4_X1   g243(.A1(G225gat), .A2(new_n417_), .A3(G233gat), .A4(new_n418_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n426_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n442_), .A2(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n416_), .A2(new_n419_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n421_), .A2(new_n426_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT95), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n428_), .A2(new_n435_), .A3(new_n420_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n434_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n433_), .A2(new_n439_), .A3(new_n447_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n457_));
  AND4_X1   g256(.A1(new_n292_), .A2(new_n299_), .A3(new_n300_), .A4(new_n456_), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n429_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n377_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n432_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n457_), .A2(new_n458_), .A3(new_n429_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n453_), .B1(new_n452_), .B2(new_n434_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n434_), .ZN(new_n465_));
  AOI211_X1 g264(.A(KEYINPUT97), .B(new_n465_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n442_), .A2(new_n443_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n446_), .A2(new_n444_), .ZN(new_n469_));
  AND4_X1   g268(.A1(new_n305_), .A2(new_n468_), .A3(new_n318_), .A4(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n463_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n471_), .A2(KEYINPUT99), .A3(new_n377_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n403_), .B1(new_n462_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT101), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT101), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n475_), .B(new_n403_), .C1(new_n462_), .C2(new_n472_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n431_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G29gat), .B(G36gat), .Z(new_n478_));
  XOR2_X1   g277(.A(G43gat), .B(G50gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n482_), .A2(KEYINPUT76), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(KEYINPUT76), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G1gat), .A2(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT14), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n483_), .A2(new_n488_), .A3(new_n486_), .A4(new_n484_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  MUX2_X1   g291(.A(new_n481_), .B(new_n480_), .S(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n492_), .B(new_n480_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n496_), .B1(new_n499_), .B2(new_n495_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT79), .ZN(new_n502_));
  XOR2_X1   g301(.A(G169gat), .B(G197gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n500_), .A2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n477_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT68), .B(G71gat), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G78gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT68), .B(G71gat), .ZN(new_n512_));
  INV_X1    g311(.A(G78gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n511_), .B(new_n514_), .C1(KEYINPUT11), .C2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT69), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n516_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n518_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n509_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G85gat), .B(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n525_), .B1(KEYINPUT9), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(KEYINPUT9), .B2(new_n525_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT6), .Z(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT10), .B(G99gat), .Z(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n525_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT7), .Z(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT67), .B(new_n537_), .C1(new_n539_), .C2(new_n532_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT8), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n521_), .A2(new_n522_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n517_), .A2(new_n518_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT70), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n524_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n536_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n530_), .A2(KEYINPUT71), .A3(new_n535_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n519_), .A2(new_n523_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT12), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n546_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT70), .B1(new_n544_), .B2(new_n545_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n542_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n547_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n562_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G176gat), .B(G204gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n571_), .B(KEYINPUT73), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT74), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n577_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n492_), .B(new_n586_), .Z(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT70), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n587_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n552_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n592_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT34), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n543_), .A2(new_n480_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n551_), .A2(new_n481_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n610_), .B(new_n609_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n613_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n616_), .B(KEYINPUT36), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT37), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n619_), .A2(new_n622_), .A3(KEYINPUT37), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n508_), .A2(new_n585_), .A3(new_n604_), .A4(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n429_), .A2(KEYINPUT102), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n429_), .A2(KEYINPUT102), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n628_), .A2(G1gat), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n477_), .A2(new_n623_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n507_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n581_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n603_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n429_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n635_), .A3(new_n641_), .ZN(G1324gat));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n636_), .A2(new_n639_), .A3(new_n643_), .A4(new_n323_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n640_), .B2(new_n322_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n322_), .A2(G8gat), .ZN(new_n650_));
  OAI22_X1  g449(.A1(new_n648_), .A2(new_n649_), .B1(new_n628_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI221_X1 g452(.A(KEYINPUT40), .B1(new_n628_), .B2(new_n650_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n640_), .B2(new_n403_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n404_), .A2(new_n397_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n628_), .B2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(new_n377_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n640_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n628_), .B2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n604_), .A2(new_n624_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT104), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n578_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n508_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n429_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n627_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n476_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT99), .B1(new_n471_), .B2(new_n377_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n455_), .A2(new_n459_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n461_), .A3(new_n660_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n675_), .A3(new_n432_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n475_), .B1(new_n676_), .B2(new_n403_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n430_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(new_n627_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n671_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n581_), .A2(new_n637_), .A3(new_n603_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n686_), .B(new_n683_), .C1(new_n671_), .C2(new_n681_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n631_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n670_), .B1(new_n688_), .B2(new_n690_), .ZN(G1328gat));
  NAND2_X1  g490(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n688_), .B2(new_n323_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n667_), .A2(new_n508_), .A3(new_n696_), .A4(new_n323_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n692_), .B(new_n695_), .C1(new_n697_), .C2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n682_), .A2(new_n684_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n686_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n323_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n698_), .B(new_n699_), .Z(new_n707_));
  NAND4_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n701_), .A2(new_n708_), .ZN(G1329gat));
  AOI21_X1  g508(.A(G43gat), .B1(new_n668_), .B2(new_n404_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n404_), .A2(G43gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n688_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g512(.A1(new_n660_), .A2(G50gat), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT108), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n668_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n688_), .A2(new_n377_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n717_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT107), .B1(new_n717_), .B2(G50gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n603_), .A2(new_n637_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n636_), .A2(new_n584_), .A3(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT109), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n724_), .B2(new_n669_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n477_), .A2(new_n637_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n581_), .A2(new_n680_), .A3(new_n603_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n728_), .A2(G57gat), .A3(new_n631_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1332gat));
  INV_X1    g529(.A(new_n728_), .ZN(new_n731_));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n323_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n724_), .A2(new_n323_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G64gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT48), .B(new_n732_), .C1(new_n724_), .C2(new_n323_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n739_), .A3(new_n404_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n724_), .A2(new_n404_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G71gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT49), .B(new_n739_), .C1(new_n724_), .C2(new_n404_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1334gat));
  NAND3_X1  g544(.A1(new_n731_), .A2(new_n513_), .A3(new_n377_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n724_), .A2(new_n377_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G78gat), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT50), .B(new_n513_), .C1(new_n724_), .C2(new_n377_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n585_), .A2(new_n666_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n726_), .ZN(new_n753_));
  INV_X1    g552(.A(G85gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n689_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n578_), .A2(new_n507_), .A3(new_n603_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT110), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n682_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n669_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n759_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g559(.A(G92gat), .B1(new_n753_), .B2(new_n323_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n323_), .A2(G92gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT111), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n758_), .B2(new_n763_), .ZN(G1337gat));
  NAND4_X1  g563(.A1(new_n752_), .A2(new_n404_), .A3(new_n534_), .A4(new_n726_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n682_), .A2(new_n757_), .A3(new_n404_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G99gat), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n767_), .A3(G99gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT51), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n766_), .B(new_n773_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n753_), .A2(new_n533_), .A3(new_n377_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n682_), .A2(new_n757_), .A3(new_n377_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1339gat));
  NAND2_X1  g582(.A1(new_n637_), .A2(new_n572_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n543_), .B1(new_n524_), .B2(new_n546_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n547_), .B(new_n553_), .C1(new_n786_), .C2(KEYINPUT12), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(new_n562_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n562_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n787_), .A2(new_n785_), .A3(new_n562_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n574_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n563_), .B1(new_n554_), .B2(new_n559_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n564_), .B1(new_n795_), .B2(new_n785_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n791_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n784_), .B1(new_n794_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n494_), .B1(new_n493_), .B2(KEYINPUT115), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(KEYINPUT115), .B2(new_n493_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n504_), .B1(new_n499_), .B2(new_n494_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n505_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT116), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n804_), .C1(new_n573_), .C2(new_n576_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n624_), .B1(new_n800_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n804_), .A2(new_n572_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n574_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n793_), .B(new_n575_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT58), .B(new_n813_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n680_), .A3(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT57), .B(new_n624_), .C1(new_n800_), .C2(new_n809_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n812_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n603_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n722_), .A2(new_n627_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n581_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n581_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n378_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n403_), .A3(new_n631_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n830_), .A2(KEYINPUT119), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n828_), .B1(new_n822_), .B2(new_n603_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n837_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n833_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT117), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(KEYINPUT59), .C1(new_n841_), .C2(new_n833_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n637_), .A2(G113gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT120), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n843_), .A2(new_n845_), .A3(new_n847_), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n830_), .A2(new_n832_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n386_), .B1(new_n851_), .B2(new_n507_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1340gat));
  NAND4_X1  g652(.A1(new_n843_), .A2(new_n845_), .A3(new_n584_), .A4(new_n847_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n841_), .A2(new_n833_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n388_), .B1(new_n581_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n856_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n388_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n603_), .A2(new_n383_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT121), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n843_), .A2(new_n845_), .A3(new_n847_), .A4(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n383_), .B1(new_n851_), .B2(new_n603_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1342gat));
  NAND4_X1  g663(.A1(new_n843_), .A2(new_n845_), .A3(new_n680_), .A4(new_n847_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G134gat), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n851_), .A2(G134gat), .A3(new_n624_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n841_), .A2(new_n404_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n323_), .A2(new_n660_), .A3(new_n631_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n507_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(G141gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n585_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n334_), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n603_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n871_), .B2(new_n627_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n623_), .A2(new_n325_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n871_), .B2(new_n881_), .ZN(G1347gat));
  AND2_X1   g681(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n841_), .A2(new_n377_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n322_), .A2(new_n403_), .A3(new_n689_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(G169gat), .B(new_n883_), .C1(new_n886_), .C2(new_n507_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n637_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT124), .Z(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n205_), .B1(new_n888_), .B2(new_n637_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n883_), .A2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n887_), .B(new_n891_), .C1(new_n892_), .C2(new_n894_), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n888_), .B2(new_n578_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n584_), .A2(G176gat), .A3(new_n885_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n896_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  NAND4_X1  g700(.A1(new_n897_), .A2(new_n898_), .A3(new_n604_), .A4(new_n885_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n603_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n902_), .A2(new_n215_), .B1(new_n888_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n886_), .B2(new_n627_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n623_), .B1(new_n231_), .B2(new_n230_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n886_), .B2(new_n906_), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n322_), .A2(new_n660_), .A3(new_n669_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n869_), .A2(new_n637_), .A3(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g709(.A1(new_n869_), .A2(new_n584_), .A3(new_n908_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n240_), .A2(KEYINPUT126), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n869_), .A2(new_n604_), .A3(new_n908_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT63), .B(G211gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n914_), .B2(new_n917_), .ZN(G1354gat));
  NAND4_X1  g717(.A1(new_n869_), .A2(new_n250_), .A3(new_n623_), .A4(new_n908_), .ZN(new_n919_));
  AND4_X1   g718(.A1(new_n403_), .A2(new_n830_), .A3(new_n680_), .A4(new_n908_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n250_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n923_), .B(new_n919_), .C1(new_n920_), .C2(new_n250_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1355gat));
endmodule


