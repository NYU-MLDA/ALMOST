//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT91), .ZN(new_n203_));
  INV_X1    g002(.A(G211gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G218gat), .ZN(new_n205_));
  INV_X1    g004(.A(G218gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G211gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(G211gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(G218gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT91), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(G204gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G197gat), .ZN(new_n215_));
  INV_X1    g014(.A(G197gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G204gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n205_), .A2(new_n207_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT90), .A4(KEYINPUT21), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n216_), .B2(G204gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n224_), .A2(KEYINPUT21), .B1(new_n215_), .B2(new_n217_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n220_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(KEYINPUT2), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n230_), .B(new_n234_), .C1(KEYINPUT2), .C2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G155gat), .B(G162gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(KEYINPUT88), .A3(new_n240_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n236_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT1), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT84), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(G155gat), .B2(G162gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(new_n249_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT85), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n248_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n243_), .A2(new_n244_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n202_), .B(new_n227_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n227_), .A2(KEYINPUT92), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT90), .B1(new_n214_), .B2(G197gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n216_), .A2(G204gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n214_), .A2(G197gat), .ZN(new_n269_));
  OAI22_X1  g068(.A1(new_n213_), .A2(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n221_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n271_), .A2(new_n220_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT92), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n266_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n243_), .A2(new_n244_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(new_n260_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n276_), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n263_), .B(new_n265_), .C1(new_n280_), .C2(new_n202_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT93), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(new_n202_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n263_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n264_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G22gat), .B(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT89), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n261_), .A2(new_n289_), .A3(new_n262_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n261_), .A2(new_n262_), .ZN(new_n297_));
  OAI211_X1 g096(.A(G228gat), .B(G233gat), .C1(new_n297_), .C2(new_n276_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n282_), .A2(new_n285_), .A3(new_n296_), .A4(new_n300_), .ZN(new_n301_));
  OAI22_X1  g100(.A1(new_n283_), .A2(new_n284_), .B1(KEYINPUT94), .B2(new_n265_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n265_), .A2(KEYINPUT94), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n263_), .A3(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n302_), .A2(new_n304_), .A3(new_n295_), .A4(new_n293_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  INV_X1    g108(.A(G176gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(KEYINPUT23), .ZN(new_n313_));
  AND2_X1   g112(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n314_));
  NOR2_X1   g113(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n312_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n311_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT26), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT25), .B(G183gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(KEYINPUT78), .A3(new_n326_), .A4(new_n328_), .ZN(new_n333_));
  INV_X1    g132(.A(G169gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n310_), .A3(KEYINPUT79), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(G169gat), .B2(G176gat), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT24), .A4(new_n307_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n316_), .A2(new_n312_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n317_), .A2(KEYINPUT23), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n335_), .A2(new_n337_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(new_n342_), .C2(KEYINPUT24), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n320_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT30), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346_));
  INV_X1    g145(.A(G43gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G15gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n345_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G113gat), .B(G120gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n354_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n306_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n344_), .A2(KEYINPUT97), .A3(new_n227_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT97), .B1(new_n344_), .B2(new_n227_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n326_), .A2(new_n328_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT95), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT95), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n332_), .A3(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n371_));
  OR2_X1    g170(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n372_));
  NAND2_X1  g171(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n317_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n312_), .A2(KEYINPUT23), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n370_), .A2(new_n376_), .A3(new_n338_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(G169gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n334_), .A2(KEYINPUT22), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT96), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n334_), .A2(KEYINPUT22), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT96), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n310_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n319_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n372_), .A2(new_n373_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n387_), .B(new_n341_), .C1(new_n388_), .C2(new_n317_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n307_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n377_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n362_), .B1(new_n365_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n344_), .A2(new_n272_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n227_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n362_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT18), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT99), .ZN(new_n403_));
  XOR2_X1   g202(.A(G64gat), .B(G92gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n400_), .A2(KEYINPUT101), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT98), .B1(new_n391_), .B2(new_n227_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n272_), .A2(new_n409_), .A3(new_n377_), .A4(new_n390_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n362_), .A2(new_n394_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OAI22_X1  g211(.A1(new_n365_), .A2(new_n412_), .B1(new_n398_), .B2(new_n397_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n407_), .B1(new_n413_), .B2(new_n406_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT101), .B1(new_n400_), .B2(new_n406_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT0), .ZN(new_n418_));
  INV_X1    g217(.A(G57gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT100), .ZN(new_n424_));
  INV_X1    g223(.A(new_n357_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n261_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n261_), .A2(new_n424_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n279_), .B2(KEYINPUT100), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n428_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n279_), .A2(new_n433_), .A3(new_n425_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n432_), .ZN(new_n437_));
  OAI221_X1 g236(.A(new_n423_), .B1(new_n430_), .B2(new_n432_), .C1(new_n435_), .C2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT102), .ZN(new_n439_));
  INV_X1    g238(.A(new_n428_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n357_), .B1(new_n261_), .B2(new_n424_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n426_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n437_), .B1(new_n442_), .B2(KEYINPUT4), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n432_), .B1(new_n434_), .B2(new_n426_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n439_), .B(new_n422_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n445_), .ZN(new_n446_));
  OAI22_X1  g245(.A1(new_n435_), .A2(new_n437_), .B1(new_n432_), .B2(new_n430_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n439_), .B1(new_n447_), .B2(new_n422_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n416_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n405_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n413_), .A2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n410_), .A2(new_n411_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n408_), .C1(new_n364_), .C2(new_n363_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n395_), .A2(new_n396_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT20), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n362_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n456_), .A3(new_n405_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n431_), .B(new_n436_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n423_), .B1(new_n442_), .B2(new_n432_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n443_), .A2(new_n444_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n423_), .ZN(new_n464_));
  NOR4_X1   g263(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT33), .A4(new_n422_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n360_), .B1(new_n449_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n359_), .B1(new_n305_), .B2(new_n301_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT27), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n413_), .A2(new_n450_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n405_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT103), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT103), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n458_), .A2(new_n474_), .A3(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n457_), .A2(KEYINPUT27), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n405_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT104), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT104), .ZN(new_n482_));
  AOI211_X1 g281(.A(new_n482_), .B(new_n479_), .C1(new_n473_), .C2(new_n475_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n468_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n359_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n306_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n446_), .A2(new_n448_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n467_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G190gat), .B(G218gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(G134gat), .B(G162gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT6), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  OR3_X1    g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(KEYINPUT8), .A3(new_n501_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT64), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n506_), .A2(KEYINPUT64), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT10), .B(G99gat), .Z(new_n510_));
  INV_X1    g309(.A(G106gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n506_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n509_), .A2(new_n512_), .A3(new_n497_), .A4(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n505_), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G29gat), .B(G36gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT34), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n521_), .B(new_n525_), .C1(new_n515_), .C2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(new_n524_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n495_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n529_), .A2(new_n494_), .A3(new_n530_), .A4(new_n493_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n531_), .B(KEYINPUT72), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n532_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n540_), .B2(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(G1gat), .ZN(new_n542_));
  INV_X1    g341(.A(G8gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G22gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G15gat), .ZN(new_n546_));
  INV_X1    g345(.A(G15gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G22gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT73), .ZN(new_n550_));
  XOR2_X1   g349(.A(G1gat), .B(G8gat), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n549_), .A2(KEYINPUT73), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(KEYINPUT73), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(KEYINPUT11), .B2(new_n560_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n559_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n569_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT74), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(new_n570_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n541_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n556_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n551_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n526_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n553_), .A2(new_n556_), .A3(new_n518_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n581_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT75), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n518_), .A2(new_n519_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n518_), .A2(new_n519_), .ZN(new_n589_));
  OAI22_X1  g388(.A1(new_n582_), .A2(new_n583_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT76), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n557_), .A2(new_n520_), .A3(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n591_), .A2(new_n581_), .A3(new_n593_), .A4(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT77), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n593_), .A2(new_n585_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n581_), .A4(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n587_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n587_), .A2(new_n598_), .A3(new_n595_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n515_), .A2(new_n567_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT66), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n567_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n611_), .A2(new_n504_), .A3(new_n505_), .A4(new_n514_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT65), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n515_), .A2(KEYINPUT66), .A3(new_n567_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n505_), .A2(new_n514_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT8), .B1(new_n500_), .B2(new_n501_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT65), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n611_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n610_), .A2(new_n613_), .A3(new_n614_), .A4(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(G230gat), .A3(G233gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n623_), .B(new_n567_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n515_), .B2(new_n567_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n622_), .B(new_n612_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT67), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n608_), .A2(KEYINPUT12), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n624_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT67), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n622_), .A4(new_n612_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n621_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G120gat), .B(G148gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT69), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n636_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n633_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n621_), .A2(new_n628_), .A3(new_n632_), .A4(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT13), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(KEYINPUT13), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR4_X1   g446(.A1(new_n490_), .A2(new_n580_), .A3(new_n607_), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n489_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n542_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n579_), .A2(new_n540_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n647_), .A2(new_n607_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT105), .B1(new_n647_), .B2(new_n607_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n306_), .A2(new_n485_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n474_), .B1(new_n458_), .B2(new_n469_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT103), .B(KEYINPUT27), .C1(new_n451_), .C2(new_n457_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n480_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n482_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n476_), .A2(KEYINPUT104), .A3(new_n480_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n661_), .A2(new_n306_), .A3(new_n485_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n489_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n467_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n657_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n489_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n651_), .A2(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n481_), .A2(new_n483_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n672_), .B(G8gat), .C1(new_n669_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n669_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n543_), .B1(new_n679_), .B2(new_n673_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n677_), .B(new_n678_), .C1(new_n672_), .C2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n648_), .A2(new_n543_), .A3(new_n673_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(KEYINPUT40), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  AOI21_X1  g486(.A(new_n547_), .B1(new_n679_), .B2(new_n485_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n689_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n648_), .A2(new_n547_), .A3(new_n485_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(G1326gat));
  OAI21_X1  g492(.A(G22gat), .B1(new_n669_), .B2(new_n306_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT42), .ZN(new_n695_));
  INV_X1    g494(.A(new_n306_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n648_), .A2(new_n545_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1327gat));
  NOR2_X1   g497(.A1(new_n579_), .A2(new_n540_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n668_), .A2(new_n653_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(G29gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n649_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n579_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n541_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(new_n541_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n668_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n703_), .B(new_n705_), .C1(new_n706_), .C2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n705_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT107), .B1(new_n711_), .B2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n668_), .B2(new_n708_), .ZN(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT43), .B(new_n541_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n704_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n703_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n710_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n649_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G29gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n718_), .B2(new_n649_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n702_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  XOR2_X1   g522(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n724_));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n718_), .B2(new_n673_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n673_), .B(KEYINPUT109), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n700_), .A2(new_n725_), .A3(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n730_));
  XOR2_X1   g529(.A(new_n729_), .B(new_n730_), .Z(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n724_), .B1(new_n726_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n724_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n674_), .B(new_n710_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n731_), .B(new_n734_), .C1(new_n735_), .C2(new_n725_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1329gat));
  AOI21_X1  g536(.A(G43gat), .B1(new_n700_), .B2(new_n485_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n359_), .A2(new_n347_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n718_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n741_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n739_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n744_), .B(new_n710_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n738_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n700_), .B2(new_n696_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n696_), .A2(G50gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n718_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n749_), .B(new_n710_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n754_), .B2(new_n748_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1331gat));
  INV_X1    g555(.A(new_n647_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n606_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n668_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n580_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n419_), .A3(new_n649_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n759_), .A2(KEYINPUT114), .A3(new_n652_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT114), .B1(new_n759_), .B2(new_n652_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n649_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n765_), .B2(new_n419_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n760_), .A2(new_n767_), .A3(new_n728_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n762_), .A2(new_n728_), .A3(new_n763_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(G64gat), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G64gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT116), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n778_), .A3(new_n485_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n764_), .A2(new_n485_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G71gat), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n760_), .A2(new_n785_), .A3(new_n696_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n764_), .A2(new_n696_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G78gat), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT50), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(KEYINPUT50), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1335gat));
  NAND2_X1  g590(.A1(new_n706_), .A2(new_n709_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n579_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n758_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT117), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n792_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n489_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n759_), .A2(new_n579_), .A3(new_n540_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n421_), .A3(new_n649_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n797_), .B2(new_n727_), .ZN(new_n802_));
  INV_X1    g601(.A(G92gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n803_), .A3(new_n673_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1337gat));
  AND3_X1   g604(.A1(new_n799_), .A2(new_n485_), .A3(new_n510_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n796_), .A2(new_n485_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(G99gat), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g608(.A1(new_n799_), .A2(new_n511_), .A3(new_n696_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n792_), .A2(new_n795_), .A3(new_n696_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  INV_X1    g616(.A(new_n581_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n591_), .A2(new_n818_), .A3(new_n593_), .A4(new_n585_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n584_), .A2(new_n585_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n604_), .B1(new_n820_), .B2(new_n581_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n605_), .A3(new_n642_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n825_), .A2(new_n605_), .A3(new_n642_), .A4(KEYINPUT121), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n627_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n622_), .B1(new_n630_), .B2(new_n612_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n628_), .A2(new_n632_), .A3(new_n831_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n639_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT56), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT122), .B1(new_n830_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n835_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n640_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n841_), .B(new_n639_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n828_), .B(new_n829_), .C1(new_n840_), .C2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n817_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n708_), .A3(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n830_), .A2(new_n837_), .A3(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n844_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT58), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n848_), .B1(new_n851_), .B2(new_n541_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n830_), .A2(new_n837_), .A3(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n643_), .A2(new_n605_), .A3(new_n825_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n840_), .A2(new_n842_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n836_), .A2(new_n856_), .A3(KEYINPUT56), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n606_), .A3(new_n642_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT57), .A3(new_n540_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n860_), .B2(new_n540_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n579_), .B1(new_n854_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n757_), .A2(new_n607_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n580_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n580_), .B2(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n649_), .B(new_n664_), .C1(new_n864_), .C2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n606_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n854_), .A2(new_n863_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n793_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n489_), .B1(new_n877_), .B2(new_n870_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n878_), .A2(KEYINPUT124), .A3(KEYINPUT59), .A4(new_n664_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n607_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n875_), .B1(new_n883_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n885_));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n647_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n873_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n757_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n886_), .ZN(G1341gat));
  INV_X1    g690(.A(G127gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n873_), .A2(new_n892_), .A3(new_n579_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n793_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n892_), .ZN(G1342gat));
  INV_X1    g694(.A(G134gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n872_), .B2(new_n540_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n899_), .B(new_n896_), .C1(new_n872_), .C2(new_n540_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n708_), .A2(G134gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1343gat));
  AND2_X1   g703(.A1(new_n727_), .A2(new_n486_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n649_), .B(new_n905_), .C1(new_n864_), .C2(new_n871_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n607_), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n907_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n757_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g709(.A1(new_n906_), .A2(new_n793_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(G162gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n906_), .B2(new_n540_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(new_n914_), .C1(new_n906_), .C2(new_n540_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n878_), .A2(G162gat), .A3(new_n708_), .A4(new_n905_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(G1347gat));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n877_), .A2(new_n870_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n727_), .A2(new_n649_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n922_), .A2(new_n468_), .A3(new_n606_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n921_), .B1(new_n925_), .B2(new_n334_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(G1348gat));
  NOR2_X1   g728(.A1(new_n864_), .A2(new_n871_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n923_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n930_), .A2(new_n658_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n647_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n579_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G183gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n332_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1350gat));
  INV_X1    g737(.A(new_n540_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n932_), .A2(new_n368_), .A3(new_n369_), .A4(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n932_), .A2(new_n708_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n942_), .B2(new_n325_), .ZN(G1351gat));
  NAND2_X1  g742(.A1(new_n923_), .A2(new_n486_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n930_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n606_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n647_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g748(.A1(new_n945_), .A2(new_n579_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n950_), .B2(new_n952_), .ZN(G1354gat));
  NAND3_X1  g752(.A1(new_n945_), .A2(G218gat), .A3(new_n708_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n944_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n922_), .A2(new_n939_), .A3(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959_));
  AOI21_X1  g758(.A(G218gat), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(KEYINPUT127), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n955_), .B1(new_n960_), .B2(new_n961_), .ZN(G1355gat));
endmodule


