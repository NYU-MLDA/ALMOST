//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G190gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT75), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G183gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n206_), .B(new_n209_), .C1(new_n212_), .C2(KEYINPUT75), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n221_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT78), .B(G169gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(G176gat), .B1(KEYINPUT77), .B2(KEYINPUT22), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n218_), .A2(new_n237_), .A3(KEYINPUT79), .A4(new_n219_), .ZN(new_n238_));
  AND2_X1   g037(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n214_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n237_), .B2(new_n217_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n236_), .B(new_n238_), .C1(new_n241_), .C2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n213_), .A2(new_n231_), .B1(new_n234_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G99gat), .ZN(new_n246_));
  INV_X1    g045(.A(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n245_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G127gat), .B(G134gat), .Z(new_n250_));
  XOR2_X1   g049(.A(G113gat), .B(G120gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n249_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(G15gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT30), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n253_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT100), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT98), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G204gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT86), .B1(new_n268_), .B2(G197gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT86), .ZN(new_n270_));
  INV_X1    g069(.A(G197gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT85), .B(G197gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n269_), .B(new_n272_), .C1(new_n273_), .C2(G204gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n267_), .B1(new_n274_), .B2(KEYINPUT21), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(KEYINPUT85), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G197gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n268_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT87), .B(new_n276_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n273_), .B2(new_n268_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT87), .B1(new_n285_), .B2(new_n276_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n275_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n285_), .A2(new_n276_), .A3(new_n266_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n218_), .A2(new_n237_), .A3(new_n219_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT79), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n227_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n292_), .A2(new_n238_), .A3(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n208_), .A2(new_n211_), .A3(new_n203_), .A4(new_n205_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n224_), .B(new_n225_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT91), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n214_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(KEYINPUT23), .B2(new_n214_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n306_), .A2(new_n236_), .B1(G169gat), .B2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT92), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n223_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n287_), .A2(new_n289_), .A3(new_n304_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT20), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n277_), .A2(new_n279_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n281_), .B1(new_n320_), .B2(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n321_), .B2(KEYINPUT21), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n282_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n288_), .B1(new_n323_), .B2(new_n275_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(new_n245_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n265_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(G204gat), .B1(new_n277_), .B2(new_n279_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n269_), .A2(new_n272_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT21), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n266_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n322_), .B2(new_n282_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n307_), .A2(new_n315_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT91), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n292_), .A2(new_n238_), .A3(new_n296_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT91), .B1(new_n298_), .B2(new_n299_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  OAI22_X1  g135(.A1(new_n331_), .A2(new_n288_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n287_), .A2(new_n245_), .A3(new_n289_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n337_), .A2(KEYINPUT20), .A3(new_n264_), .A4(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G8gat), .B(G36gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n261_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  AOI211_X1 g145(.A(KEYINPUT98), .B(new_n344_), .C1(new_n326_), .C2(new_n339_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT27), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n333_), .A2(new_n335_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n349_), .A2(new_n297_), .B1(new_n307_), .B2(new_n315_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n338_), .B(KEYINPUT20), .C1(new_n324_), .C2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n265_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n324_), .B2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n287_), .A2(new_n289_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n245_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n264_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n352_), .A2(new_n344_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT99), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n352_), .A2(new_n358_), .A3(KEYINPUT99), .A4(new_n344_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n260_), .B1(new_n348_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n351_), .A2(new_n265_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n264_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n345_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT98), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n340_), .A2(new_n261_), .A3(new_n345_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n362_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(KEYINPUT100), .A3(KEYINPUT27), .A4(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n344_), .B1(new_n352_), .B2(new_n358_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT27), .B1(new_n375_), .B2(new_n359_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT81), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n386_), .A2(new_n388_), .B1(new_n384_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT80), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n396_), .A2(KEYINPUT3), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(KEYINPUT81), .A3(new_n385_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n390_), .A2(new_n395_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n405_), .A2(new_n401_), .A3(KEYINPUT83), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n396_), .A2(new_n387_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n401_), .B1(KEYINPUT1), .B2(new_n403_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n403_), .A2(KEYINPUT1), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n413_), .A3(new_n252_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT94), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n399_), .B2(new_n407_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(new_n252_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n416_), .A2(KEYINPUT94), .A3(new_n252_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n383_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n416_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n252_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n416_), .B2(new_n252_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n419_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT95), .A3(new_n383_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n425_), .A2(KEYINPUT4), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n383_), .B(new_n433_), .C1(new_n430_), .C2(KEYINPUT4), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n382_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(KEYINPUT4), .ZN(new_n436_));
  INV_X1    g235(.A(new_n383_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n433_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(new_n381_), .A3(new_n422_), .A4(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G22gat), .B(G50gat), .Z(new_n442_));
  NOR3_X1   g241(.A1(new_n423_), .A2(KEYINPUT29), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n416_), .B2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n416_), .A2(new_n445_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n324_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n448_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n355_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n450_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n443_), .A2(new_n446_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n449_), .B1(new_n324_), .B2(new_n448_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G228gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(G78gat), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n454_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n441_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n373_), .A2(new_n377_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n352_), .A2(new_n358_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n340_), .B2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n441_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n440_), .A2(KEYINPUT96), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n432_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(KEYINPUT96), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n381_), .A3(new_n439_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484_));
  INV_X1    g283(.A(new_n359_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(new_n374_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n375_), .A2(KEYINPUT93), .A3(new_n359_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n383_), .B1(new_n430_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n488_), .B2(new_n430_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n436_), .A2(new_n383_), .A3(new_n438_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n382_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n477_), .B1(new_n483_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n470_), .A2(new_n466_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n259_), .B1(new_n472_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n372_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT27), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT100), .B1(new_n500_), .B2(new_n371_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n495_), .B(new_n377_), .C1(new_n498_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT101), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n376_), .B1(new_n364_), .B2(new_n372_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n495_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n259_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n441_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n497_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT71), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519_));
  INV_X1    g318(.A(G1gat), .ZN(new_n520_));
  INV_X1    g319(.A(G8gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n517_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n517_), .B(new_n525_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G113gat), .B(G141gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n534_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n510_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT7), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT6), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT8), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT67), .B1(new_n545_), .B2(new_n550_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT8), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n548_), .B(KEYINPUT66), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n541_), .B(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(KEYINPUT68), .B2(new_n544_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n544_), .A2(KEYINPUT68), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI22_X1  g360(.A1(new_n553_), .A2(new_n554_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n551_), .B(new_n552_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n561_), .A2(new_n555_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(KEYINPUT69), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT10), .B(G99gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT64), .ZN(new_n570_));
  INV_X1    g369(.A(G106gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n546_), .B1(new_n573_), .B2(new_n547_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n547_), .A2(new_n573_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT65), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT65), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n579_), .A3(new_n544_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n568_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(KEYINPUT12), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n562_), .A2(new_n580_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT12), .B1(new_n591_), .B2(new_n589_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n580_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n594_), .B2(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n589_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT5), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT70), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n597_), .A2(new_n601_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n605_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT70), .A3(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT13), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n612_), .A3(KEYINPUT13), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n517_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT72), .B1(new_n591_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n594_), .A2(new_n620_), .A3(new_n517_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n593_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n518_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n619_), .B(new_n621_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT35), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n624_), .A2(new_n625_), .B1(KEYINPUT36), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n624_), .B2(KEYINPUT73), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n619_), .A2(new_n621_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n581_), .A2(new_n518_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT73), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .A4(new_n632_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n629_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n628_), .A2(KEYINPUT36), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n629_), .A2(new_n634_), .A3(new_n639_), .A4(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n642_), .A2(KEYINPUT37), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT37), .B1(new_n642_), .B2(new_n644_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n525_), .B(new_n588_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT17), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G127gat), .B(G155gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT16), .ZN(new_n654_));
  XOR2_X1   g453(.A(G183gat), .B(G211gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(KEYINPUT17), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT74), .Z(new_n660_));
  NOR2_X1   g459(.A1(new_n648_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n540_), .A2(new_n617_), .A3(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT102), .Z(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n441_), .A2(new_n520_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n642_), .A2(new_n644_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n510_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT105), .ZN(new_n672_));
  INV_X1    g471(.A(new_n660_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n617_), .A2(new_n538_), .A3(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT104), .Z(new_n675_));
  AND3_X1   g474(.A1(new_n672_), .A2(KEYINPUT106), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT106), .B1(new_n672_), .B2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n441_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n666_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n668_), .A2(new_n680_), .A3(new_n681_), .ZN(G1324gat));
  INV_X1    g481(.A(new_n504_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n521_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n683_), .A3(new_n675_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G8gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G8gat), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n665_), .A2(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI221_X1 g490(.A(KEYINPUT40), .B1(new_n687_), .B2(new_n688_), .C1(new_n665_), .C2(new_n684_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n678_), .B2(new_n508_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n663_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT107), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n696_), .A3(new_n698_), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n495_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n663_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G22gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G22gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n617_), .A2(new_n538_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n510_), .B2(new_n647_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(new_n509_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n648_), .B(new_n710_), .C1(new_n712_), .C2(new_n497_), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n673_), .B(new_n708_), .C1(new_n709_), .C2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(KEYINPUT44), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(G29gat), .A3(new_n441_), .ZN(new_n719_));
  INV_X1    g518(.A(G29gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n669_), .A2(new_n673_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n540_), .A2(new_n617_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n679_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n719_), .A2(new_n723_), .ZN(G1328gat));
  NOR3_X1   g523(.A1(new_n722_), .A2(G36gat), .A3(new_n504_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n716_), .A2(new_n683_), .A3(new_n717_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G36gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n728_), .B(new_n729_), .Z(G1329gat));
  NOR2_X1   g529(.A1(new_n508_), .A2(new_n247_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n717_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n716_), .A2(KEYINPUT110), .A3(new_n717_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n247_), .B1(new_n722_), .B2(new_n508_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT47), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1330gat));
  NAND3_X1  g542(.A1(new_n718_), .A2(G50gat), .A3(new_n701_), .ZN(new_n744_));
  INV_X1    g543(.A(G50gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n722_), .B2(new_n495_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1331gat));
  NOR2_X1   g546(.A1(new_n617_), .A2(new_n538_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n510_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n661_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n679_), .B1(new_n751_), .B2(KEYINPUT112), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(KEYINPUT112), .B2(new_n751_), .ZN(new_n753_));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n672_), .A2(new_n673_), .A3(new_n748_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n679_), .A2(new_n754_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT113), .Z(G1332gat));
  INV_X1    g557(.A(G64gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n755_), .B2(new_n683_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n683_), .A2(new_n759_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n762_), .A2(new_n763_), .B1(new_n751_), .B2(new_n764_), .ZN(G1333gat));
  NAND2_X1  g564(.A1(new_n755_), .A2(new_n259_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G71gat), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT49), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n508_), .A2(G71gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n751_), .B2(new_n769_), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n755_), .A2(new_n701_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G78gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT50), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n495_), .A2(G78gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n751_), .B2(new_n774_), .ZN(G1335gat));
  AND2_X1   g574(.A1(new_n750_), .A2(new_n721_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n441_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n617_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n539_), .A3(new_n660_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n709_), .B2(new_n713_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n441_), .A2(G85gat), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT115), .Z(new_n782_));
  AOI21_X1  g581(.A(new_n777_), .B1(new_n780_), .B2(new_n782_), .ZN(G1336gat));
  AOI21_X1  g582(.A(G92gat), .B1(new_n776_), .B2(new_n683_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n683_), .A2(G92gat), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT116), .Z(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n780_), .B2(new_n786_), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n776_), .A2(new_n259_), .A3(new_n570_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n780_), .A2(new_n259_), .ZN(new_n789_));
  INV_X1    g588(.A(G99gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g591(.A1(new_n776_), .A2(new_n571_), .A3(new_n701_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n495_), .B(new_n779_), .C1(new_n709_), .C2(new_n713_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n571_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n779_), .ZN(new_n798_));
  AND4_X1   g597(.A1(new_n505_), .A2(new_n373_), .A3(new_n377_), .A4(new_n495_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n505_), .B1(new_n504_), .B2(new_n495_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n509_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n472_), .A2(new_n496_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n508_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n710_), .B1(new_n804_), .B2(new_n648_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT43), .B(new_n647_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n701_), .B(new_n798_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n794_), .B1(new_n797_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G106gat), .B1(new_n807_), .B2(KEYINPUT117), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n796_), .B1(new_n780_), .B2(new_n701_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(KEYINPUT52), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n793_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT119), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n810_), .B2(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n780_), .A2(new_n796_), .A3(new_n701_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n808_), .A2(new_n816_), .A3(new_n794_), .A4(G106gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n793_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n821_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n818_), .B2(new_n793_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n793_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT119), .B(new_n825_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n822_), .A2(new_n827_), .ZN(G1339gat));
  AOI21_X1  g627(.A(new_n596_), .B1(new_n590_), .B2(new_n595_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n597_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n590_), .A2(new_n595_), .A3(KEYINPUT55), .A4(new_n596_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n606_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(KEYINPUT120), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n607_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n538_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n534_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n527_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n537_), .B1(new_n531_), .B2(new_n529_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n841_), .A2(new_n537_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n610_), .A2(new_n612_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n669_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n835_), .A2(new_n844_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n837_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n647_), .B1(new_n850_), .B2(KEYINPUT58), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n848_), .B(new_n852_), .C1(new_n849_), .C2(new_n837_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n846_), .A2(new_n847_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n669_), .C1(new_n840_), .C2(new_n845_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n673_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n661_), .A2(new_n539_), .A3(new_n617_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n507_), .A2(new_n441_), .A3(new_n259_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT122), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n538_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(KEYINPUT59), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n539_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n871_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873_));
  AOI21_X1  g672(.A(G120gat), .B1(new_n778_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(G120gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n865_), .B(new_n875_), .C1(new_n874_), .C2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n617_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n865_), .A2(new_n882_), .A3(new_n673_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n660_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n882_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n865_), .B2(new_n670_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n868_), .A2(new_n870_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT124), .B(G134gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n647_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n887_), .B2(new_n889_), .ZN(G1343gat));
  NAND4_X1  g689(.A1(new_n504_), .A2(new_n701_), .A3(new_n441_), .A4(new_n508_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n860_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n860_), .A2(new_n894_), .A3(new_n891_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n538_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g696(.A(new_n778_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g698(.A(new_n673_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  NOR2_X1   g701(.A1(new_n893_), .A2(new_n895_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G162gat), .B1(new_n903_), .B2(new_n647_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n669_), .A2(G162gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(new_n905_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n854_), .A2(new_n855_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n660_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n857_), .B(KEYINPUT54), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n504_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n701_), .A2(new_n711_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n314_), .A3(new_n538_), .A4(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n683_), .B(new_n911_), .C1(new_n856_), .C2(new_n859_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G169gat), .B1(new_n913_), .B2(new_n539_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n914_), .A3(KEYINPUT62), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(new_n919_), .C1(KEYINPUT62), .C2(new_n914_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n913_), .A2(new_n617_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT127), .B(G176gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n922_), .B(new_n923_), .Z(G1349gat));
  NOR2_X1   g723(.A1(new_n913_), .A2(new_n660_), .ZN(new_n925_));
  MUX2_X1   g724(.A(G183gat), .B(new_n212_), .S(new_n925_), .Z(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n913_), .B2(new_n647_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n670_), .A2(new_n206_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n913_), .B2(new_n928_), .ZN(G1351gat));
  NAND3_X1  g728(.A1(new_n910_), .A2(new_n508_), .A3(new_n471_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n539_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n271_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n617_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n268_), .ZN(G1353gat));
  NAND2_X1  g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n673_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n930_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n930_), .B2(new_n647_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n669_), .A2(G218gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n930_), .B2(new_n941_), .ZN(G1355gat));
endmodule


