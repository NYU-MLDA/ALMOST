//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(G71gat), .ZN(new_n203_));
  INV_X1    g002(.A(G78gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT71), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT71), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G71gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n209_), .A3(new_n204_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G78gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n203_), .A2(new_n204_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT11), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n216_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT11), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G1gat), .A2(G8gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT14), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G1gat), .ZN(new_n225_));
  INV_X1    g024(.A(G8gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n222_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n221_), .A2(new_n222_), .A3(new_n227_), .A4(new_n223_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n220_), .B(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(G231gat), .A2(G233gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G155gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT16), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G211gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT76), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n240_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT6), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT6), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G99gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT10), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT10), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G99gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT65), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n249_), .A2(new_n251_), .A3(KEYINPUT68), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G85gat), .ZN(new_n270_));
  INV_X1    g069(.A(G92gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n269_), .A2(new_n272_), .A3(KEYINPUT67), .A4(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n254_), .A2(new_n265_), .A3(new_n266_), .A4(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n267_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n277_), .B(KEYINPUT9), .C1(new_n276_), .C2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT69), .B1(new_n275_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n266_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT68), .B1(new_n249_), .B2(new_n251_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n278_), .A2(new_n276_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n285_), .A2(new_n273_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .A4(new_n279_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n272_), .A2(new_n267_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT8), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n254_), .A2(new_n266_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n291_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n296_), .A2(new_n298_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(KEYINPUT70), .A3(new_n295_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n290_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT8), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n297_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G43gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G29gat), .A2(G36gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G43gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G29gat), .A2(G36gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n305_), .A2(G50gat), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(G50gat), .B1(new_n305_), .B2(new_n310_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n289_), .A2(new_n303_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n310_), .ZN(new_n315_));
  INV_X1    g114(.A(G50gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n305_), .A2(G50gat), .A3(new_n310_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT15), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT15), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n289_), .A2(new_n303_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n314_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n296_), .A2(new_n298_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n252_), .A3(new_n300_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n290_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT8), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n328_), .A2(new_n297_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT72), .B1(new_n329_), .B2(new_n313_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n323_), .A2(new_n331_), .A3(KEYINPUT73), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G232gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT34), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT35), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n323_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(KEYINPUT35), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n289_), .A2(new_n303_), .A3(new_n313_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n321_), .A2(new_n319_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n329_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n330_), .B1(KEYINPUT72), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n337_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n343_), .B(KEYINPUT73), .C1(new_n344_), .C2(new_n335_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G190gat), .B(G218gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G134gat), .ZN(new_n348_));
  INV_X1    g147(.A(G162gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT36), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT74), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n350_), .B(KEYINPUT36), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n338_), .A2(new_n345_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n352_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT37), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT37), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n338_), .A2(new_n345_), .A3(new_n355_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n364_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n356_), .A2(KEYINPUT75), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n247_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT77), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G120gat), .B(G148gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT5), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G176gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G230gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT64), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n329_), .A2(new_n220_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n289_), .A2(new_n303_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n220_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n381_), .A3(KEYINPUT12), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n220_), .B1(new_n289_), .B2(new_n303_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT12), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n377_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n377_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n375_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n289_), .A2(new_n303_), .A3(new_n220_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n390_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n385_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n375_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n389_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT13), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT13), .B1(new_n389_), .B2(new_n396_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n231_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n340_), .B2(new_n231_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G229gat), .A2(G233gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n231_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n321_), .B2(new_n319_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n405_), .ZN(new_n409_));
  NOR4_X1   g208(.A1(new_n408_), .A2(KEYINPUT78), .A3(new_n403_), .A4(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n313_), .A2(new_n407_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n413_), .B2(new_n403_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G141gat), .ZN(new_n415_));
  INV_X1    g214(.A(G169gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G197gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .A4(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n311_), .A2(new_n312_), .A3(new_n320_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT15), .B1(new_n317_), .B2(new_n318_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n231_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n403_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n405_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT78), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n404_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n414_), .A4(new_n418_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT80), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n419_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n418_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n401_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT3), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n442_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT2), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  OR2_X1    g247(.A1(G155gat), .A2(G162gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n448_), .A2(KEYINPUT1), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(KEYINPUT1), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n437_), .A2(new_n438_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n444_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G120gat), .ZN(new_n457_));
  INV_X1    g256(.A(G127gat), .ZN(new_n458_));
  INV_X1    g257(.A(G134gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G113gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G127gat), .A2(G134gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n457_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G120gat), .A3(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n456_), .A2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n450_), .A2(new_n468_), .A3(new_n466_), .A4(new_n455_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT94), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n450_), .A2(new_n455_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474_));
  INV_X1    g273(.A(new_n469_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n470_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n472_), .A2(new_n478_), .A3(new_n476_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n482_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT18), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G64gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(new_n271_), .ZN(new_n495_));
  AND2_X1   g294(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n237_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n500_), .A2(KEYINPUT91), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT91), .B1(new_n500_), .B2(new_n501_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(G169gat), .B2(G176gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G176gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT24), .B1(new_n416_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT92), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n416_), .A3(new_n509_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(new_n511_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G183gat), .A2(G190gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n514_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n505_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n504_), .A2(new_n515_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n416_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(G169gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT93), .ZN(new_n530_));
  INV_X1    g329(.A(G190gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n237_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n518_), .A2(new_n519_), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n528_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G197gat), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G211gat), .B(G218gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537_));
  OR3_X1    g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G197gat), .B(G204gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT21), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n537_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n536_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n524_), .A2(new_n534_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n533_), .A2(KEYINPUT83), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT83), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n518_), .A2(new_n532_), .A3(new_n545_), .A4(new_n519_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n529_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT25), .B1(new_n237_), .B2(KEYINPUT81), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT81), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n499_), .A3(G183gat), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n548_), .B(new_n550_), .C1(new_n497_), .C2(new_n496_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n506_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n523_), .A2(new_n551_), .A3(new_n552_), .A4(new_n520_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n538_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G226gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT19), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR4_X1   g359(.A1(new_n543_), .A2(new_n556_), .A3(new_n557_), .A4(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n524_), .A2(new_n538_), .A3(new_n542_), .A4(new_n534_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n495_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n494_), .B(G92gat), .ZN(new_n566_));
  NOR4_X1   g365(.A1(new_n543_), .A2(new_n556_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n569_), .A3(KEYINPUT27), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571_));
  INV_X1    g370(.A(new_n564_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n524_), .A2(new_n534_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n555_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n556_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(KEYINPUT20), .A4(new_n559_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n566_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n565_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT27), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n571_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI211_X1 g379(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n565_), .C2(new_n577_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n491_), .B(new_n570_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT84), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n547_), .A2(new_n553_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n554_), .A2(KEYINPUT84), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n547_), .A2(new_n553_), .A3(new_n585_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(KEYINPUT30), .A3(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n588_), .A2(new_n591_), .A3(KEYINPUT86), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT86), .B1(new_n588_), .B2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G227gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n206_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G15gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT85), .B(G99gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G43gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n596_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n592_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n588_), .A2(new_n591_), .A3(KEYINPUT86), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT87), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n469_), .B(KEYINPUT31), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n593_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT87), .ZN(new_n609_));
  INV_X1    g408(.A(new_n603_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT87), .B(new_n605_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G78gat), .B(G106gat), .ZN(new_n614_));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT29), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n555_), .B1(new_n473_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT89), .B(G233gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G228gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(KEYINPUT90), .A3(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(KEYINPUT90), .Z(new_n623_));
  OAI211_X1 g422(.A(new_n555_), .B(new_n623_), .C1(new_n473_), .C2(new_n618_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n617_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n456_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT28), .B1(new_n456_), .B2(KEYINPUT29), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G50gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n316_), .A3(new_n628_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n624_), .A3(new_n617_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n626_), .A2(new_n630_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n631_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(new_n625_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n612_), .A2(new_n613_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n583_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT32), .B(new_n495_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n561_), .A2(new_n564_), .B1(new_n566_), .B2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n641_), .B(new_n643_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n482_), .A2(new_n488_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n487_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(KEYINPUT33), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n490_), .A2(KEYINPUT96), .A3(KEYINPUT33), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n477_), .A2(new_n481_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n478_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n472_), .A2(new_n476_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n653_), .B(new_n487_), .C1(new_n654_), .C2(new_n478_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n578_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n655_), .B(new_n656_), .C1(new_n490_), .C2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n644_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n633_), .A2(new_n636_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n613_), .B2(new_n612_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n435_), .B1(new_n640_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n370_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n491_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n225_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT38), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n435_), .B(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n640_), .A2(new_n662_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n366_), .A2(new_n367_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n247_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n670_), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n491_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT100), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n667_), .A2(new_n676_), .ZN(G1324gat));
  OR2_X1    g476(.A1(new_n580_), .A2(new_n581_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n570_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n664_), .A2(new_n226_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G8gat), .B1(new_n674_), .B2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(KEYINPUT39), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(KEYINPUT39), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT101), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n680_), .B(new_n687_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  NAND2_X1  g490(.A1(new_n612_), .A2(new_n613_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G15gat), .B1(new_n674_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT41), .Z(new_n694_));
  INV_X1    g493(.A(G15gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n692_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n664_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT102), .Z(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n674_), .B2(new_n637_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n664_), .A2(new_n615_), .A3(new_n660_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n671_), .A2(new_n246_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n663_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n665_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n669_), .A2(new_n247_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n709_));
  AOI21_X1  g508(.A(new_n359_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT74), .B(new_n357_), .C1(new_n338_), .C2(new_n345_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n363_), .B1(new_n712_), .B2(new_n356_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n353_), .A2(KEYINPUT75), .A3(new_n356_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n367_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT37), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT104), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n362_), .A2(new_n368_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n709_), .B1(new_n720_), .B2(new_n670_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n713_), .A2(new_n716_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(KEYINPUT105), .A3(new_n723_), .A4(new_n670_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n670_), .A2(new_n362_), .A3(new_n723_), .A4(new_n368_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n708_), .B1(new_n721_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n708_), .B(KEYINPUT44), .C1(new_n721_), .C2(new_n728_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n665_), .A2(G29gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n707_), .B1(new_n733_), .B2(new_n734_), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n679_), .A3(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT106), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n731_), .A2(new_n738_), .A3(new_n679_), .A4(new_n732_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(G36gat), .A3(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n679_), .B(KEYINPUT107), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n705_), .A2(G36gat), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT45), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n740_), .A2(KEYINPUT46), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1329gat));
  OAI21_X1  g547(.A(new_n308_), .B1(new_n705_), .B2(new_n692_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n731_), .A2(G43gat), .A3(new_n696_), .A4(new_n732_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n750_), .A2(new_n751_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n755_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(new_n316_), .B1(new_n733_), .B2(new_n660_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n705_), .A2(G50gat), .A3(new_n637_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n760_), .A2(KEYINPUT110), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT110), .B1(new_n760_), .B2(new_n761_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1331gat));
  INV_X1    g563(.A(new_n401_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n434_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n670_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n370_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n665_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771_));
  INV_X1    g570(.A(new_n673_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n767_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n768_), .A2(KEYINPUT111), .A3(new_n673_), .ZN(new_n774_));
  AND4_X1   g573(.A1(G57gat), .A2(new_n773_), .A3(new_n665_), .A4(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n770_), .A2(new_n775_), .ZN(G1332gat));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n741_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n778_), .A3(new_n774_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G64gat), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n206_), .A3(new_n696_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n773_), .A2(new_n696_), .A3(new_n774_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G71gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n786_), .A3(G71gat), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(KEYINPUT49), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT49), .B1(new_n789_), .B2(new_n790_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n785_), .B1(new_n791_), .B2(new_n792_), .ZN(G1334gat));
  NAND3_X1  g592(.A1(new_n769_), .A2(new_n204_), .A3(new_n660_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n773_), .A2(new_n660_), .A3(new_n774_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G78gat), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT50), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT50), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1335gat));
  NAND2_X1  g598(.A1(new_n768_), .A2(new_n704_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n665_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n721_), .A2(new_n728_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n246_), .A2(new_n401_), .A3(new_n434_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n491_), .A2(new_n270_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(G1336gat));
  AOI21_X1  g607(.A(G92gat), .B1(new_n801_), .B2(new_n679_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n741_), .A2(new_n271_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n806_), .B2(new_n810_), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n805_), .B2(new_n692_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n259_), .A3(new_n696_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n803_), .A2(new_n660_), .A3(new_n804_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G106gat), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n801_), .A2(new_n264_), .A3(new_n660_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n819_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n816_), .A2(G106gat), .A3(new_n822_), .A4(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n821_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT53), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n820_), .A2(new_n827_), .A3(new_n821_), .A4(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n393_), .A2(KEYINPUT55), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n386_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n391_), .A2(new_n392_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n830_), .A2(new_n832_), .B1(new_n377_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n395_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n377_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n386_), .A2(new_n831_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT55), .B(new_n377_), .C1(new_n382_), .C2(new_n385_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n375_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n835_), .A2(new_n396_), .A3(new_n841_), .A4(new_n434_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n422_), .A2(KEYINPUT115), .A3(new_n423_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n408_), .B2(new_n403_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n845_), .A3(new_n409_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n418_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n405_), .B1(new_n413_), .B2(new_n403_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n419_), .B2(new_n428_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n397_), .A2(new_n850_), .A3(KEYINPUT116), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n397_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n842_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n671_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n395_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n840_), .B1(new_n839_), .B2(new_n375_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT58), .A3(new_n396_), .A4(new_n850_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n835_), .A2(new_n396_), .A3(new_n841_), .A4(new_n850_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n862_), .A2(new_n368_), .A3(new_n362_), .A4(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n855_), .A2(KEYINPUT57), .A3(new_n671_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n858_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n247_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n434_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n246_), .B(new_n870_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT114), .B1(new_n871_), .B2(KEYINPUT54), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(KEYINPUT54), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n369_), .A2(new_n874_), .A3(new_n875_), .A4(new_n870_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n873_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n869_), .A2(new_n877_), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n679_), .A2(new_n491_), .A3(new_n692_), .A4(new_n660_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT59), .ZN(new_n881_));
  INV_X1    g680(.A(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n858_), .A2(new_n866_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT117), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n858_), .A2(new_n866_), .A3(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n867_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n882_), .B1(new_n887_), .B2(new_n247_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n879_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n881_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n891_), .A2(new_n461_), .A3(new_n766_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n434_), .A3(new_n879_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n461_), .B2(new_n893_), .ZN(G1340gat));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n858_), .A2(new_n866_), .A3(new_n885_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n885_), .B1(new_n858_), .B2(new_n866_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n867_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n877_), .B1(new_n899_), .B2(new_n246_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n890_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n900_), .A2(new_n901_), .B1(KEYINPUT59), .B2(new_n880_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n457_), .B1(new_n902_), .B2(new_n765_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n457_), .A2(KEYINPUT60), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT60), .B1(new_n765_), .B2(new_n457_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n880_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n895_), .B1(new_n903_), .B2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G120gat), .B1(new_n891_), .B2(new_n401_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n906_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(KEYINPUT118), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1341gat));
  OAI21_X1  g710(.A(G127gat), .B1(new_n891_), .B2(new_n247_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n882_), .A2(new_n246_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n879_), .A2(new_n458_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1342gat));
  INV_X1    g714(.A(new_n722_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n891_), .A2(new_n459_), .A3(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n878_), .A2(new_n672_), .A3(new_n879_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n459_), .B2(new_n918_), .ZN(G1343gat));
  NAND3_X1  g718(.A1(new_n741_), .A2(new_n665_), .A3(new_n639_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT119), .Z(new_n921_));
  NAND2_X1  g720(.A1(new_n878_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n766_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT120), .B(G141gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1344gat));
  NOR2_X1   g724(.A1(new_n922_), .A2(new_n401_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT121), .B(G148gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1345gat));
  NAND3_X1  g727(.A1(new_n882_), .A2(new_n921_), .A3(new_n246_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  OAI21_X1  g730(.A(new_n349_), .B1(new_n922_), .B2(new_n671_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n878_), .A2(G162gat), .A3(new_n720_), .A4(new_n921_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT122), .ZN(G1347gat));
  INV_X1    g734(.A(KEYINPUT22), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n741_), .A2(new_n665_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n638_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n900_), .A2(new_n936_), .A3(new_n434_), .A4(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(G169gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n888_), .A2(new_n766_), .A3(new_n938_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n941_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n416_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n942_), .B2(new_n946_), .ZN(G1348gat));
  NAND4_X1  g746(.A1(new_n878_), .A2(new_n939_), .A3(G176gat), .A4(new_n765_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n888_), .A2(new_n401_), .A3(new_n938_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(G176gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR2_X1   g750(.A1(new_n913_), .A2(new_n938_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n953_), .B1(new_n237_), .B2(new_n952_), .ZN(G1350gat));
  NAND4_X1  g753(.A1(new_n900_), .A2(new_n498_), .A3(new_n672_), .A4(new_n939_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n888_), .A2(new_n916_), .A3(new_n938_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n531_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT125), .ZN(G1351gat));
  AND2_X1   g757(.A1(new_n937_), .A2(new_n639_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n960_), .B1(new_n869_), .B2(new_n877_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(new_n434_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n765_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n374_), .A2(KEYINPUT126), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n964_), .B(new_n965_), .ZN(G1353gat));
  NOR2_X1   g765(.A1(new_n913_), .A2(new_n960_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n967_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968_));
  XOR2_X1   g767(.A(KEYINPUT63), .B(G211gat), .Z(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n967_), .B2(new_n969_), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n961_), .B2(new_n672_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n722_), .A2(G218gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n961_), .B2(new_n972_), .ZN(new_n973_));
  XOR2_X1   g772(.A(new_n973_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


