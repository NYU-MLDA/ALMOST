//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G231gat), .ZN(new_n210_));
  INV_X1    g009(.A(G233gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  XOR2_X1   g013(.A(G71gat), .B(G78gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n214_), .A2(new_n215_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n219_), .B(new_n212_), .C1(new_n217_), .C2(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT73), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n219_), .B1(new_n217_), .B2(new_n216_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n226_), .B2(new_n221_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n209_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT73), .B1(new_n220_), .B2(new_n222_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n224_), .A3(new_n221_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n208_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G155gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G183gat), .B(G211gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n241_), .A3(new_n239_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT17), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n228_), .A2(new_n247_), .A3(new_n232_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n251_), .A2(KEYINPUT6), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(KEYINPUT6), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT10), .B(G99gat), .Z(new_n255_));
  INV_X1    g054(.A(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G85gat), .A2(G92gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT9), .ZN(new_n259_));
  OR2_X1    g058(.A1(G85gat), .A2(G92gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(KEYINPUT9), .A3(new_n258_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n254_), .A2(new_n257_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(G85gat), .A2(G92gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G85gat), .A2(G92gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT64), .B1(new_n260_), .B2(new_n258_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  OR3_X1    g068(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n268_), .A2(new_n269_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n269_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n262_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT65), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT15), .ZN(new_n277_));
  XOR2_X1   g076(.A(G29gat), .B(G36gat), .Z(new_n278_));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G29gat), .B(G36gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT70), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n277_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT15), .A3(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n262_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n276_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT34), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT35), .ZN(new_n296_));
  AND4_X1   g095(.A1(new_n254_), .A2(new_n257_), .A3(new_n261_), .A4(new_n259_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n268_), .A2(new_n272_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT8), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n268_), .A2(new_n269_), .A3(new_n272_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n285_), .A2(new_n286_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n296_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(KEYINPUT35), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT69), .Z(new_n305_));
  AND3_X1   g104(.A1(new_n293_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n293_), .B2(new_n303_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G190gat), .B(G218gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT36), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT71), .Z(new_n313_));
  NOR3_X1   g112(.A1(new_n306_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n310_), .B(KEYINPUT36), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT72), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n321_), .B(new_n317_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n314_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n323_), .B2(KEYINPUT37), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n250_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n225_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT12), .B1(new_n275_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT66), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(KEYINPUT12), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n276_), .A3(new_n292_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n301_), .A2(new_n225_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n275_), .A2(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G176gat), .B(G204gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT68), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n336_), .A2(new_n340_), .A3(new_n347_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT13), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT13), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n353_), .A3(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n326_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(KEYINPUT76), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n208_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G229gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n302_), .B2(new_n208_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n302_), .B(new_n208_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n361_), .A2(new_n364_), .B1(new_n365_), .B2(new_n363_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(KEYINPUT77), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G141gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G169gat), .B(G197gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n367_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT81), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT30), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n380_), .B(new_n381_), .C1(new_n384_), .C2(KEYINPUT24), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT79), .B(G190gat), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n389_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n389_), .B2(KEYINPUT26), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT78), .B(G183gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n393_), .ZN(new_n397_));
  INV_X1    g196(.A(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(KEYINPUT26), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n388_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n389_), .A2(new_n396_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n402_));
  OAI21_X1  g201(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(G71gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n407_), .A2(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n377_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n376_), .A3(new_n413_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G134gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G127gat), .ZN(new_n422_));
  INV_X1    g221(.A(G127gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G134gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G120gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G113gat), .ZN(new_n427_));
  INV_X1    g226(.A(G113gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G120gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n422_), .A2(new_n424_), .A3(new_n427_), .A4(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT83), .ZN(new_n439_));
  INV_X1    g238(.A(new_n431_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT31), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n420_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n416_), .A2(new_n418_), .A3(KEYINPUT85), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n420_), .B2(new_n446_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT18), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  AND2_X1   g255(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(G197gat), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G197gat), .A2(G204gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT21), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G211gat), .B(G218gat), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT90), .B(G204gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n460_), .B1(new_n466_), .B2(G197gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT91), .B1(new_n467_), .B2(KEYINPUT21), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n469_), .A3(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n464_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n466_), .A2(G197gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n463_), .B1(G197gat), .B2(G204gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n465_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT96), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n405_), .A2(new_n478_), .A3(new_n403_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n394_), .A2(new_n398_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n380_), .A2(new_n381_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n405_), .B2(new_n403_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n477_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(KEYINPUT97), .A3(new_n481_), .A4(new_n479_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT24), .B1(new_n382_), .B2(new_n383_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n487_), .A2(KEYINPUT95), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n487_), .A2(KEYINPUT95), .B1(new_n382_), .B2(new_n383_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n385_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT25), .B(G183gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G190gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT94), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n491_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n484_), .A2(new_n486_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT98), .B1(new_n476_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n469_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT91), .B(KEYINPUT21), .C1(new_n459_), .C2(new_n461_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n475_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n465_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n484_), .A2(new_n486_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n490_), .A2(new_n498_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n407_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n466_), .A2(G197gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n474_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n464_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n465_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT92), .B1(new_n503_), .B2(new_n504_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n511_), .A2(new_n520_), .A3(KEYINPUT20), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G226gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT19), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n517_), .B1(new_n516_), .B2(new_n465_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n503_), .A2(KEYINPUT92), .A3(new_n504_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n407_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT20), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n476_), .B2(new_n499_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n456_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n526_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n512_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n528_), .B1(new_n535_), .B2(new_n511_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n456_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n452_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n452_), .B1(new_n541_), .B2(new_n456_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n482_), .A2(new_n483_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n498_), .B2(new_n490_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n533_), .B1(new_n476_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n527_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n523_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n511_), .A2(new_n520_), .A3(KEYINPUT20), .A4(new_n528_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n546_), .B2(new_n523_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n537_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n542_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(G155gat), .A2(G162gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G155gat), .A2(G162gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT88), .B1(new_n559_), .B2(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(G141gat), .A2(G148gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT3), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G141gat), .A2(G148gat), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT2), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n564_), .A2(new_n567_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n561_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n562_), .B2(new_n572_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT87), .B1(new_n557_), .B2(KEYINPUT1), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT1), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(G155gat), .A4(G162gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n557_), .A2(KEYINPUT1), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n576_), .A2(new_n579_), .A3(new_n555_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n571_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT29), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n505_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(G228gat), .A3(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G228gat), .A2(G233gat), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n525_), .A2(new_n526_), .A3(new_n584_), .A4(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G22gat), .B(G50gat), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n561_), .A2(new_n570_), .B1(new_n575_), .B2(new_n581_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT28), .B1(new_n583_), .B2(KEYINPUT29), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n591_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G78gat), .B(G106gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(KEYINPUT93), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n586_), .B(new_n590_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n597_), .A2(new_n601_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n586_), .A2(new_n590_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n437_), .A2(new_n442_), .A3(new_n583_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n431_), .A2(new_n432_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n592_), .A2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n616_), .A2(KEYINPUT4), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT4), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n437_), .A2(new_n442_), .A3(new_n620_), .A4(new_n583_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G225gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n615_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G1gat), .B(G29gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT100), .B(G85gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT0), .B(G57gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n616_), .A2(new_n618_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n622_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n616_), .A2(KEYINPUT4), .A3(new_n618_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n634_), .A2(KEYINPUT99), .A3(new_n623_), .A4(new_n621_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n625_), .A2(new_n631_), .A3(new_n633_), .A4(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n625_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n630_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n614_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n540_), .A2(new_n553_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n636_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n541_), .A2(new_n641_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n630_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n625_), .A2(new_n633_), .A3(new_n635_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n632_), .A2(new_n623_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n634_), .A2(new_n622_), .A3(new_n621_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n630_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n524_), .A2(new_n456_), .A3(new_n531_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n537_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n636_), .A2(new_n647_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .A4(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n614_), .B1(new_n646_), .B2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n451_), .B1(new_n640_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n451_), .A2(new_n644_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n540_), .A2(new_n553_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n614_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n373_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n358_), .A2(KEYINPUT76), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n359_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n644_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(G1gat), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT103), .Z(new_n672_));
  XOR2_X1   g471(.A(new_n323_), .B(KEYINPUT104), .Z(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n372_), .A2(new_n675_), .A3(new_n250_), .A4(new_n355_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n203_), .B1(new_n676_), .B2(new_n644_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n672_), .A2(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(new_n661_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n204_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT39), .Z(new_n682_));
  INV_X1    g481(.A(new_n666_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n204_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n451_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n676_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT105), .Z(G1326gat));
  INV_X1    g492(.A(G22gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n676_), .B2(new_n614_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT42), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n683_), .A2(new_n694_), .A3(new_n614_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1327gat));
  NOR3_X1   g497(.A1(new_n356_), .A2(new_n250_), .A3(new_n373_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n324_), .B2(KEYINPUT106), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n325_), .B(new_n701_), .C1(new_n659_), .C2(new_n663_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n659_), .A2(new_n663_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n324_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n699_), .B1(new_n702_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n699_), .C1(new_n702_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n667_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n323_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n356_), .A2(new_n712_), .A3(new_n250_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n664_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n714_), .A2(G29gat), .A3(new_n667_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n711_), .A2(new_n715_), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n714_), .A2(G36gat), .A3(new_n661_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT45), .Z(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n708_), .A2(new_n719_), .A3(new_n680_), .A4(new_n709_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n708_), .A2(new_n680_), .A3(new_n709_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT107), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  AND4_X1   g523(.A1(KEYINPUT108), .A2(new_n723_), .A3(G36gat), .A4(new_n720_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n718_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n718_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND2_X1  g529(.A1(new_n688_), .A2(G43gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n714_), .A2(new_n451_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n710_), .A2(new_n731_), .B1(G43gat), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g533(.A(G50gat), .B1(new_n710_), .B2(new_n662_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n662_), .A2(G50gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT109), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n714_), .B2(new_n737_), .ZN(G1331gat));
  AOI21_X1  g537(.A(new_n372_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n325_), .A2(new_n739_), .A3(new_n250_), .A4(new_n356_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n644_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n675_), .A2(new_n373_), .A3(new_n250_), .A4(new_n356_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT110), .Z(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n644_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n742_), .B1(new_n745_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n744_), .B2(new_n680_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n747_), .A3(new_n680_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1333gat));
  AOI21_X1  g550(.A(new_n409_), .B1(new_n744_), .B2(new_n688_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT49), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n740_), .A2(new_n409_), .A3(new_n688_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n744_), .B2(new_n614_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n740_), .A2(new_n756_), .A3(new_n614_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1335gat));
  INV_X1    g560(.A(new_n250_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n739_), .A2(new_n323_), .A3(new_n762_), .A4(new_n356_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT112), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n644_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n702_), .A2(new_n705_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n373_), .A3(new_n356_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n644_), .A2(G85gat), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT114), .Z(new_n771_));
  AOI21_X1  g570(.A(new_n766_), .B1(new_n769_), .B2(new_n771_), .ZN(G1336gat));
  INV_X1    g571(.A(G92gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n764_), .A2(new_n773_), .A3(new_n680_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n767_), .A2(new_n661_), .A3(new_n768_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n773_), .ZN(G1337gat));
  AND3_X1   g575(.A1(new_n764_), .A2(new_n688_), .A3(new_n255_), .ZN(new_n777_));
  INV_X1    g576(.A(G99gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n769_), .B2(new_n688_), .ZN(new_n779_));
  OAI22_X1  g578(.A1(new_n777_), .A2(new_n779_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n780_));
  NAND2_X1  g579(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1338gat));
  AND3_X1   g581(.A1(new_n764_), .A2(new_n256_), .A3(new_n614_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n769_), .A2(new_n614_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT116), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n769_), .A2(new_n786_), .A3(new_n614_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(G106gat), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT52), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n785_), .A2(new_n790_), .A3(G106gat), .A4(new_n787_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n783_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n793_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n783_), .B(new_n795_), .C1(new_n789_), .C2(new_n791_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  AND3_X1   g596(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n373_), .B1(new_n798_), .B2(new_n245_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n325_), .B(new_n355_), .C1(new_n799_), .C2(KEYINPUT118), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n250_), .B2(new_n373_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT54), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n356_), .A2(new_n324_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n799_), .A2(KEYINPUT118), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n250_), .A2(new_n801_), .A3(new_n373_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT12), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n337_), .A2(KEYINPUT66), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n328_), .A2(KEYINPUT66), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n333_), .B(new_n332_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n810_), .B1(new_n815_), .B2(new_n339_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n339_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n815_), .A2(new_n810_), .A3(new_n339_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n348_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT56), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n335_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n336_), .B1(new_n822_), .B2(new_n810_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n347_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n821_), .A2(new_n827_), .A3(new_n372_), .A4(new_n350_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n365_), .A2(new_n362_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n371_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n362_), .B1(new_n302_), .B2(new_n208_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n830_), .A2(KEYINPUT119), .B1(new_n361_), .B2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n831_), .A2(new_n833_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n351_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n712_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n350_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n840_));
  AOI211_X1 g639(.A(KEYINPUT56), .B(new_n347_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(KEYINPUT58), .A4(new_n834_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n821_), .A2(new_n827_), .A3(new_n350_), .A4(new_n834_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT120), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n325_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n844_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n836_), .A2(KEYINPUT57), .A3(new_n712_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n839_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n809_), .B1(new_n851_), .B2(new_n762_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n667_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n680_), .A2(new_n614_), .A3(new_n451_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n428_), .A3(new_n372_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n373_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n857_), .B1(new_n861_), .B2(new_n428_), .ZN(G1340gat));
  OAI21_X1  g661(.A(new_n426_), .B1(new_n355_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n856_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n426_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n355_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n426_), .ZN(G1341gat));
  OAI21_X1  g665(.A(new_n423_), .B1(new_n855_), .B2(new_n762_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n868_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n858_), .A2(new_n860_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n250_), .A2(G127gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT122), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n856_), .A2(new_n421_), .A3(new_n674_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n325_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n421_), .ZN(G1343gat));
  NOR3_X1   g676(.A1(new_n680_), .A2(new_n662_), .A3(new_n688_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n853_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n372_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n356_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n879_), .A2(new_n762_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  AOI21_X1  g686(.A(G162gat), .B1(new_n880_), .B2(new_n674_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n324_), .A2(G162gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT123), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n880_), .B2(new_n890_), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n851_), .A2(new_n762_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n809_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n661_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n660_), .A2(new_n662_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n836_), .B2(new_n712_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n838_), .B(new_n323_), .C1(new_n828_), .C2(new_n835_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n250_), .B1(new_n901_), .B2(new_n849_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n680_), .B(new_n897_), .C1(new_n902_), .C2(new_n809_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n898_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT22), .B(G169gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n372_), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n903_), .B2(new_n373_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT124), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n911_), .B(G169gat), .C1(new_n903_), .C2(new_n373_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n909_), .A2(new_n910_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n907_), .B1(new_n913_), .B2(new_n914_), .ZN(G1348gat));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n383_), .A3(new_n356_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G176gat), .B1(new_n903_), .B2(new_n355_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1349gat));
  NOR2_X1   g717(.A1(new_n762_), .A2(new_n491_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n894_), .A2(new_n250_), .A3(new_n897_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n905_), .A2(new_n919_), .B1(new_n396_), .B2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(new_n674_), .B1(new_n497_), .B2(new_n494_), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT126), .Z(new_n923_));
  AOI21_X1  g722(.A(new_n895_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n852_), .A2(KEYINPUT125), .A3(new_n661_), .A4(new_n896_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n325_), .B1(new_n898_), .B2(new_n904_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n398_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT127), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n926_), .B(new_n930_), .C1(new_n927_), .C2(new_n398_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n894_), .A2(new_n639_), .A3(new_n451_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n372_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n933_), .A2(new_n355_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(G204gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n466_), .B2(new_n937_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(new_n933_), .A2(new_n762_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1354gat));
  OR3_X1    g742(.A1(new_n933_), .A2(G218gat), .A3(new_n673_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G218gat), .B1(new_n933_), .B2(new_n325_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1355gat));
endmodule


