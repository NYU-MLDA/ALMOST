//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT99), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT27), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G226gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT19), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT94), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT75), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT76), .B(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n207_), .B1(new_n219_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(KEYINPUT94), .A3(new_n218_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  MUX2_X1   g035(.A(new_n235_), .B(KEYINPUT24), .S(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n211_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n213_), .A2(new_n214_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(KEYINPUT23), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n227_), .A2(new_n229_), .B1(new_n234_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G204gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n247_), .B2(G204gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G211gat), .B(G218gat), .Z(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT21), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n256_), .A4(new_n251_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n247_), .B2(G204gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n245_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n248_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n253_), .B1(new_n261_), .B2(KEYINPUT21), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(new_n246_), .A3(new_n256_), .A4(new_n248_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT87), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n257_), .A2(new_n262_), .A3(new_n268_), .A4(new_n265_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n255_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n244_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n242_), .A2(new_n210_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n223_), .A3(new_n222_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n233_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT26), .B(G190gat), .Z(new_n275_));
  OAI221_X1 g074(.A(new_n237_), .B1(new_n274_), .B2(new_n275_), .C1(new_n217_), .C2(new_n215_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n206_), .B1(new_n271_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n267_), .A2(new_n269_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n254_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(new_n277_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n206_), .B1(new_n244_), .B2(new_n270_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G8gat), .B(G36gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n280_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n280_), .B2(new_n286_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n204_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n227_), .A2(new_n229_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n234_), .A2(new_n243_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n281_), .B1(new_n283_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n206_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n270_), .A2(new_n278_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n228_), .A2(new_n218_), .ZN(new_n302_));
  AND4_X1   g101(.A1(new_n282_), .A2(new_n254_), .A3(new_n296_), .A4(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n278_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n206_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n291_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n280_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT27), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT82), .ZN(new_n314_));
  INV_X1    g113(.A(G141gat), .ZN(new_n315_));
  INV_X1    g114(.A(G148gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT3), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n314_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n319_), .ZN(new_n326_));
  AND3_X1   g125(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n321_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT82), .ZN(new_n329_));
  OR2_X1    g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n325_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n331_), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT81), .B1(new_n331_), .B2(KEYINPUT1), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(KEYINPUT1), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .A4(new_n330_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G134gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G127gat), .ZN(new_n343_));
  INV_X1    g142(.A(G127gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G134gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G120gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G113gat), .ZN(new_n348_));
  INV_X1    g147(.A(G113gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G120gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(KEYINPUT78), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT78), .B1(new_n352_), .B2(new_n353_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n341_), .A2(new_n357_), .ZN(new_n358_));
  AND4_X1   g157(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n343_), .A2(new_n345_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT96), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT96), .B1(new_n359_), .B2(new_n360_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n334_), .A2(new_n361_), .A3(new_n340_), .A4(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n313_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT4), .B1(new_n341_), .B2(new_n357_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n312_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n311_), .A3(new_n363_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G85gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT0), .B(G57gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n367_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n371_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n366_), .A2(KEYINPUT98), .A3(new_n367_), .A4(new_n371_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n294_), .A2(new_n310_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT77), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT31), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n354_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n386_), .B2(new_n354_), .ZN(new_n389_));
  OAI21_X1  g188(.A(G99gat), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(G71gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT31), .B1(new_n355_), .B2(new_n356_), .ZN(new_n394_));
  INV_X1    g193(.A(G99gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n387_), .A3(new_n354_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n390_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n390_), .B2(new_n397_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n384_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n277_), .B(KEYINPUT79), .Z(new_n401_));
  INV_X1    g200(.A(new_n393_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n388_), .A2(new_n389_), .A3(G99gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n390_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n384_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n400_), .A2(new_n401_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n401_), .B1(new_n400_), .B2(new_n408_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n381_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n401_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n398_), .A2(new_n399_), .A3(new_n384_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n407_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n400_), .A2(new_n401_), .A3(new_n408_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT80), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G228gat), .ZN(new_n418_));
  INV_X1    g217(.A(G233gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n326_), .A2(new_n328_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n332_), .B1(new_n422_), .B2(new_n314_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n423_), .A2(new_n329_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n341_), .A2(KEYINPUT89), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n420_), .B1(new_n429_), .B2(new_n270_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT90), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n420_), .B1(new_n341_), .B2(KEYINPUT29), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n283_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G22gat), .B(G50gat), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n424_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n424_), .B2(new_n438_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n435_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n431_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n430_), .A2(new_n434_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n430_), .A2(KEYINPUT91), .A3(new_n434_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n432_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n420_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT89), .B1(new_n341_), .B2(new_n427_), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n421_), .B(new_n425_), .C1(new_n334_), .C2(new_n340_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n459_), .B2(new_n283_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n434_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n455_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n447_), .B1(new_n462_), .B2(new_n435_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n411_), .B(new_n417_), .C1(new_n454_), .C2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n409_), .A2(new_n410_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n444_), .A2(new_n446_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n283_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n467_), .A2(new_n420_), .B1(new_n283_), .B2(new_n433_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(new_n432_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n431_), .B1(new_n468_), .B2(KEYINPUT91), .ZN(new_n470_));
  INV_X1    g269(.A(new_n453_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(new_n435_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n466_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n380_), .B1(new_n464_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n372_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n311_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n358_), .A2(new_n363_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT97), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n312_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n480_), .A2(new_n481_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n376_), .B(new_n479_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT33), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n478_), .B1(new_n486_), .B2(new_n372_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n292_), .A2(new_n293_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n280_), .A2(new_n286_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n487_), .A2(new_n488_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n411_), .A2(new_n472_), .A3(new_n417_), .A4(new_n474_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n476_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT72), .B(G15gat), .ZN(new_n500_));
  INV_X1    g299(.A(G22gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G1gat), .A2(G8gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT14), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G29gat), .B(G36gat), .Z(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n506_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n499_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n510_), .B(KEYINPUT15), .ZN(new_n516_));
  INV_X1    g315(.A(new_n511_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n505_), .A2(new_n506_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n512_), .A3(new_n498_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G113gat), .B(G141gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT74), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G169gat), .B(G197gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n203_), .B1(new_n497_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT99), .B(new_n531_), .C1(new_n476_), .C2(new_n496_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT37), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n508_), .B(new_n509_), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT15), .ZN(new_n537_));
  XOR2_X1   g336(.A(G85gat), .B(G92gat), .Z(new_n538_));
  NOR2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n538_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT8), .ZN(new_n546_));
  INV_X1    g345(.A(new_n544_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  INV_X1    g347(.A(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n538_), .A2(KEYINPUT9), .ZN(new_n551_));
  INV_X1    g350(.A(G85gat), .ZN(new_n552_));
  INV_X1    g351(.A(G92gat), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT9), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n547_), .A2(new_n550_), .A3(new_n551_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n546_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n537_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n536_), .B(new_n555_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n557_), .A2(KEYINPUT69), .A3(new_n562_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n555_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n569_), .B2(new_n563_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n566_), .B(new_n562_), .C1(new_n570_), .C2(new_n516_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n557_), .A2(new_n566_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n560_), .B(KEYINPUT35), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n567_), .A2(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n567_), .A2(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n574_), .A2(new_n575_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT70), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n576_), .A2(KEYINPUT70), .A3(new_n585_), .ZN(new_n588_));
  AOI221_X4 g387(.A(new_n535_), .B1(new_n577_), .B2(new_n581_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n577_), .A2(new_n581_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n534_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT67), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT64), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT11), .ZN(new_n598_));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n597_), .A2(KEYINPUT11), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n596_), .B1(new_n556_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT65), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n556_), .A2(new_n605_), .A3(new_n603_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n603_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT65), .B1(new_n570_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n570_), .A2(KEYINPUT64), .A3(new_n607_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n604_), .A2(new_n606_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n570_), .B2(new_n607_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n556_), .B2(new_n603_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n607_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G120gat), .B(G148gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n613_), .A2(new_n618_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n595_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT67), .B(KEYINPUT13), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n625_), .A3(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G127gat), .B(G155gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT16), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT17), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n603_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n507_), .A2(new_n511_), .A3(new_n607_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n642_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n641_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n647_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(new_n645_), .A3(new_n640_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT73), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n649_), .A2(new_n645_), .B1(new_n640_), .B2(new_n639_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT73), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n646_), .A2(new_n647_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n652_), .B(new_n653_), .C1(new_n654_), .C2(new_n640_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n593_), .A2(new_n633_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n533_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT100), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n533_), .A2(new_n660_), .A3(new_n657_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n379_), .A2(G1gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT101), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n663_), .A2(KEYINPUT101), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n202_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT38), .A3(new_n664_), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n529_), .B(new_n656_), .C1(new_n628_), .C2(new_n632_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n584_), .A2(new_n586_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n585_), .B1(new_n576_), .B2(KEYINPUT70), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n591_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n670_), .B(new_n674_), .C1(new_n476_), .C2(new_n496_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n379_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n667_), .A2(new_n669_), .A3(new_n676_), .ZN(G1324gat));
  XNOR2_X1  g476(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n310_), .A2(new_n294_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G8gat), .B1(new_n675_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT102), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(G8gat), .C1(new_n675_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n688_), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n681_), .A2(G8gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n659_), .A2(new_n661_), .A3(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n690_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n691_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n679_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n690_), .A2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT104), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n678_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1325gat));
  NAND2_X1  g500(.A1(new_n411_), .A2(new_n417_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G15gat), .B1(new_n675_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT41), .Z(new_n705_));
  AND2_X1   g504(.A1(new_n659_), .A2(new_n661_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n703_), .A2(G15gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n450_), .A2(new_n451_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n431_), .A3(new_n453_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n711_), .A2(new_n469_), .B1(new_n473_), .B2(new_n466_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G22gat), .B1(new_n675_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n501_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n707_), .B2(new_n717_), .ZN(G1327gat));
  NAND2_X1  g517(.A1(new_n673_), .A2(new_n656_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n633_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n533_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G29gat), .B1(new_n721_), .B2(new_n493_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n656_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n633_), .A2(new_n529_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n475_), .B1(new_n702_), .B2(new_n712_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n380_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n487_), .A2(new_n488_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n492_), .A2(new_n493_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n712_), .A3(new_n703_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n725_), .B1(new_n733_), .B2(new_n593_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n593_), .B(new_n725_), .C1(new_n476_), .C2(new_n496_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n724_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT44), .B(new_n724_), .C1(new_n734_), .C2(new_n736_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n493_), .A2(G29gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n722_), .B1(new_n741_), .B2(new_n742_), .ZN(G1328gat));
  NOR2_X1   g542(.A1(new_n681_), .A2(G36gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT99), .B1(new_n733_), .B2(new_n531_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n532_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n720_), .B(new_n744_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT107), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n533_), .A2(new_n749_), .A3(new_n720_), .A4(new_n744_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n748_), .A2(KEYINPUT45), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n748_), .B2(new_n750_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n680_), .A3(new_n740_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n754_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT106), .B1(new_n754_), .B2(G36gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI221_X1 g558(.A(new_n753_), .B1(KEYINPUT108), .B2(KEYINPUT46), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1329gat));
  NAND2_X1  g560(.A1(new_n739_), .A2(new_n740_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n465_), .A2(G43gat), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n721_), .A2(new_n702_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n762_), .A2(new_n763_), .B1(new_n764_), .B2(G43gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(G1330gat));
  AOI21_X1  g566(.A(G50gat), .B1(new_n721_), .B2(new_n716_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n716_), .A2(G50gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n741_), .B2(new_n769_), .ZN(G1331gat));
  NOR2_X1   g569(.A1(new_n497_), .A2(new_n531_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n593_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n633_), .A3(new_n723_), .A4(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G57gat), .B1(new_n774_), .B2(new_n493_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n497_), .A2(new_n673_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n633_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n651_), .A2(new_n655_), .A3(new_n529_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G57gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n493_), .B2(KEYINPUT110), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(KEYINPUT110), .B2(new_n782_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n775_), .B1(new_n781_), .B2(new_n784_), .ZN(G1332gat));
  OAI21_X1  g584(.A(G64gat), .B1(new_n780_), .B2(new_n681_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT48), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n681_), .A2(G64gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n773_), .B2(new_n788_), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n780_), .B2(new_n703_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT49), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n774_), .A2(new_n392_), .A3(new_n702_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1334gat));
  OAI21_X1  g592(.A(G78gat), .B1(new_n780_), .B2(new_n712_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT50), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n712_), .A2(G78gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n773_), .B2(new_n796_), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n734_), .A2(new_n736_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n723_), .A2(new_n531_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n633_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802_), .B2(new_n379_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n771_), .A2(new_n633_), .A3(new_n656_), .A4(new_n673_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n552_), .A3(new_n493_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1336gat));
  OAI21_X1  g606(.A(G92gat), .B1(new_n802_), .B2(new_n681_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n553_), .A3(new_n680_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n802_), .B2(new_n703_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n465_), .A3(new_n548_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(KEYINPUT111), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n813_), .B(new_n815_), .ZN(G1338gat));
  NAND3_X1  g615(.A1(new_n805_), .A2(new_n549_), .A3(new_n716_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n549_), .B1(new_n801_), .B2(new_n716_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n817_), .B(new_n823_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT54), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n778_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n673_), .A2(new_n535_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n590_), .A2(new_n591_), .A3(new_n534_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n830_), .A2(KEYINPUT113), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n633_), .B2(new_n778_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n828_), .A2(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n833_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n829_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n616_), .A2(new_n617_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n604_), .A2(new_n609_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n612_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n618_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT55), .B(new_n614_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n623_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT56), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n850_), .A3(new_n623_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n498_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n519_), .A2(new_n512_), .A3(new_n499_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n524_), .A3(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n625_), .A2(new_n526_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n851_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n849_), .A2(KEYINPUT58), .A3(new_n851_), .A4(new_n855_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n593_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n848_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n626_), .A2(new_n529_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n847_), .A2(KEYINPUT115), .A3(new_n850_), .A4(new_n623_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n862_), .A2(new_n849_), .A3(new_n863_), .A4(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n526_), .B(new_n854_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n673_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n860_), .B1(new_n867_), .B2(KEYINPUT57), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n867_), .A2(KEYINPUT57), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n656_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n840_), .A2(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n475_), .A2(new_n680_), .A3(new_n379_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n349_), .A3(new_n531_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(KEYINPUT59), .A3(new_n872_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n872_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n876_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n873_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT116), .A3(new_n877_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n529_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n875_), .B1(new_n884_), .B2(new_n349_), .ZN(G1340gat));
  OAI21_X1  g684(.A(new_n347_), .B1(new_n777_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n874_), .B(new_n886_), .C1(KEYINPUT60), .C2(new_n347_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n777_), .B1(new_n882_), .B2(new_n877_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n347_), .ZN(G1341gat));
  NAND3_X1  g688(.A1(new_n874_), .A2(new_n344_), .A3(new_n723_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n656_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n344_), .ZN(G1342gat));
  NAND3_X1  g691(.A1(new_n874_), .A2(new_n342_), .A3(new_n673_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n772_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n342_), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n464_), .A2(new_n379_), .A3(new_n680_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT117), .Z(new_n897_));
  NAND2_X1  g696(.A1(new_n871_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n529_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n315_), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n777_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n316_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n656_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  INV_X1    g704(.A(G162gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n898_), .A2(new_n906_), .A3(new_n772_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n898_), .B2(new_n674_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n908_), .A2(KEYINPUT118), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(KEYINPUT118), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n909_), .B2(new_n910_), .ZN(G1347gat));
  NAND2_X1  g710(.A1(new_n680_), .A2(new_n379_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n912_), .A2(new_n703_), .A3(new_n716_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n871_), .A2(KEYINPUT119), .A3(new_n531_), .A4(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G169gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n913_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n840_), .B2(new_n870_), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT119), .B1(new_n917_), .B2(new_n531_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n915_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n871_), .A2(new_n531_), .A3(new_n913_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n922_), .A2(new_n923_), .A3(G169gat), .A4(new_n914_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n919_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT121), .B(new_n925_), .C1(new_n915_), .C2(new_n918_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n871_), .A2(new_n913_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT122), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n917_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n933_), .A2(new_n221_), .A3(new_n531_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n927_), .A2(new_n928_), .A3(new_n934_), .ZN(G1348gat));
  AND3_X1   g734(.A1(new_n917_), .A2(G176gat), .A3(new_n633_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n936_), .A2(KEYINPUT123), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(KEYINPUT123), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n933_), .A2(new_n633_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n937_), .A2(new_n938_), .B1(new_n939_), .B2(new_n220_), .ZN(G1349gat));
  AOI21_X1  g739(.A(G183gat), .B1(new_n917_), .B2(new_n723_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n933_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n723_), .A2(new_n274_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT124), .B(new_n942_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n930_), .B2(new_n932_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n941_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n945_), .A2(new_n948_), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n943_), .B2(new_n772_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n933_), .A2(new_n232_), .A3(new_n673_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n912_), .A2(new_n464_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n871_), .A2(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n529_), .ZN(new_n955_));
  OR2_X1    g754(.A1(new_n247_), .A2(KEYINPUT125), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n247_), .A2(KEYINPUT125), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n955_), .B2(new_n957_), .ZN(G1352gat));
  NOR2_X1   g758(.A1(new_n954_), .A2(new_n777_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT126), .B(G204gat), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1353gat));
  INV_X1    g761(.A(new_n954_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964_));
  INV_X1    g763(.A(G211gat), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n723_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(KEYINPUT127), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n963_), .A2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n964_), .A2(new_n965_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n968_), .B(new_n969_), .ZN(G1354gat));
  OR3_X1    g769(.A1(new_n954_), .A2(G218gat), .A3(new_n674_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G218gat), .B1(new_n954_), .B2(new_n772_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1355gat));
endmodule


