//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215_));
  NOR4_X1   g014(.A1(KEYINPUT87), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n215_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G141gat), .ZN(new_n226_));
  INV_X1    g025(.A(G148gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT3), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n218_), .A2(new_n219_), .A3(new_n217_), .ZN(new_n230_));
  AND4_X1   g029(.A1(new_n215_), .A2(new_n229_), .A3(new_n224_), .A4(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n211_), .B(new_n214_), .C1(new_n225_), .C2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT1), .B1(new_n208_), .B2(new_n209_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n209_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n207_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n214_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n218_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G127gat), .A2(G134gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G127gat), .A2(G134gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G113gat), .ZN(new_n244_));
  INV_X1    g043(.A(G113gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(G120gat), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(G120gat), .B1(new_n244_), .B2(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n232_), .A2(new_n240_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT97), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n232_), .A2(new_n240_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n254_), .A2(KEYINPUT97), .A3(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT4), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT98), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n214_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n229_), .A2(new_n224_), .A3(new_n230_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT88), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n229_), .A2(new_n224_), .A3(new_n215_), .A4(new_n230_), .ZN(new_n268_));
  AOI211_X1 g067(.A(new_n210_), .B(new_n265_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n240_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n255_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n232_), .A2(new_n240_), .A3(new_n249_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT97), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n265_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n211_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n252_), .A3(new_n249_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n260_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n206_), .B1(new_n264_), .B2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n262_), .B1(new_n277_), .B2(KEYINPUT4), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n273_), .A2(new_n276_), .B1(G225gat), .B2(G233gat), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n205_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT79), .A3(new_n285_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n288_), .A2(KEYINPUT24), .A3(new_n292_), .A4(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT25), .B(G183gat), .ZN(new_n297_));
  INV_X1    g096(.A(G190gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT77), .B1(new_n298_), .B2(KEYINPUT26), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n297_), .B(new_n299_), .C1(new_n300_), .C2(KEYINPUT77), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305_));
  INV_X1    g104(.A(new_n295_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT79), .B1(new_n294_), .B2(new_n285_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT81), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT82), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(KEYINPUT23), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n311_), .A2(new_n317_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n308_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n296_), .A2(KEYINPUT80), .A3(new_n301_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n304_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(KEYINPUT23), .A3(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n309_), .A2(new_n312_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n290_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n332_), .A3(new_n292_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT30), .ZN(new_n335_));
  XOR2_X1   g134(.A(G71gat), .B(G99gat), .Z(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n335_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n249_), .B(KEYINPUT31), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT84), .B1(new_n345_), .B2(KEYINPUT83), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(KEYINPUT84), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n283_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT95), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  OR2_X1    g158(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n329_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n290_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT94), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n363_), .A2(new_n292_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n291_), .A2(KEYINPUT94), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n288_), .A2(new_n292_), .A3(new_n295_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n297_), .A2(new_n300_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n325_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n364_), .A2(new_n365_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G197gat), .ZN(new_n375_));
  INV_X1    g174(.A(G197gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G204gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(KEYINPUT91), .B2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n375_), .A2(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(KEYINPUT90), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n378_), .A2(new_n384_), .A3(KEYINPUT21), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT21), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n375_), .B(new_n377_), .C1(KEYINPUT90), .C2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n373_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n357_), .B1(new_n372_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n334_), .A2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT19), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n319_), .A2(new_n327_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT95), .B1(new_n330_), .B2(new_n331_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n360_), .A2(new_n359_), .A3(new_n329_), .ZN(new_n398_));
  AOI21_X1  g197(.A(G176gat), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n292_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n401_), .A3(new_n365_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n368_), .A2(new_n325_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n357_), .B1(new_n404_), .B2(new_n389_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n395_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n322_), .A2(new_n333_), .A3(new_n390_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n393_), .A2(new_n395_), .B1(new_n408_), .B2(KEYINPUT100), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT20), .B1(new_n404_), .B2(new_n389_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n390_), .B1(new_n322_), .B2(new_n333_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT100), .B(new_n395_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n356_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n405_), .A2(new_n407_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n395_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n391_), .A2(new_n392_), .A3(new_n406_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n355_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(KEYINPUT27), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT102), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n410_), .A2(new_n411_), .A3(new_n395_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n356_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n418_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI211_X1 g225(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n423_), .C2(new_n418_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n419_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G22gat), .B(G50gat), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n275_), .B2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n254_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n275_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT28), .B1(new_n254_), .B2(KEYINPUT29), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n430_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n390_), .B2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n389_), .C1(new_n275_), .C2(new_n433_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n389_), .A2(KEYINPUT89), .B1(G228gat), .B2(G233gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n433_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n390_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G78gat), .B(G106gat), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  NOR4_X1   g251(.A1(new_n440_), .A2(new_n450_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n437_), .A2(new_n438_), .A3(new_n430_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n452_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n451_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n456_), .A2(new_n458_), .B1(new_n459_), .B2(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n453_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n429_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n350_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n348_), .A2(new_n349_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n257_), .A2(new_n467_), .A3(new_n260_), .A4(new_n259_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n206_), .B1(new_n277_), .B2(new_n261_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n258_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n259_), .A2(new_n260_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT99), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n278_), .B(new_n206_), .C1(new_n470_), .C2(new_n262_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n423_), .A2(new_n418_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n264_), .A2(KEYINPUT33), .A3(new_n278_), .A4(new_n206_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n416_), .A2(new_n417_), .A3(new_n480_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n482_), .B(new_n483_), .C1(new_n279_), .C2(new_n282_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n462_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT101), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT102), .B1(new_n477_), .B2(KEYINPUT27), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n424_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n205_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n450_), .A2(KEYINPUT92), .ZN(new_n492_));
  OAI22_X1  g291(.A1(new_n492_), .A2(new_n440_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n456_), .A2(KEYINPUT92), .A3(new_n459_), .A4(new_n457_), .ZN(new_n494_));
  AND4_X1   g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n474_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT103), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n490_), .A2(new_n495_), .A3(new_n496_), .A4(new_n419_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n461_), .A2(new_n283_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT103), .B1(new_n428_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT101), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n485_), .A2(new_n500_), .A3(new_n462_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n487_), .A2(new_n497_), .A3(new_n499_), .A4(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n464_), .B1(new_n466_), .B2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G57gat), .B(G64gat), .Z(new_n504_));
  INV_X1    g303(.A(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(G71gat), .A2(G78gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT67), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n504_), .A2(new_n505_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n509_), .A2(KEYINPUT67), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(KEYINPUT67), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G85gat), .B(G92gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT6), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n520_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n522_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT10), .B(G99gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  INV_X1    g334(.A(G92gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(KEYINPUT9), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT64), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT64), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n534_), .B(new_n540_), .C1(KEYINPUT9), .C2(new_n537_), .ZN(new_n541_));
  AOI211_X1 g340(.A(new_n531_), .B(new_n533_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n530_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n517_), .A2(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n513_), .B(new_n516_), .C1(new_n530_), .C2(new_n542_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT12), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n531_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(G106gat), .B2(new_n532_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n528_), .B(KEYINPUT8), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n516_), .A4(new_n513_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n544_), .A2(new_n545_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n374_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n290_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT13), .B1(new_n564_), .B2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G29gat), .B(G36gat), .ZN(new_n571_));
  INV_X1    g370(.A(G43gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G50gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G15gat), .B(G22gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G1gat), .A2(G8gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT14), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G1gat), .B(G8gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G50gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n573_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT15), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT15), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n574_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n582_), .B1(new_n588_), .B2(new_n581_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n574_), .A2(new_n581_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT75), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT76), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT74), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n245_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n598_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n570_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n517_), .B(new_n580_), .ZN(new_n611_));
  AND2_X1   g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(KEYINPUT17), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT72), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n613_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT73), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n619_), .B(KEYINPUT17), .Z(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n620_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n503_), .A2(new_n610_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G134gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G162gat), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(KEYINPUT36), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n588_), .A2(new_n550_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n548_), .A2(new_n549_), .A3(new_n584_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT68), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT34), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(KEYINPUT35), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n633_), .A2(new_n640_), .A3(new_n641_), .A4(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n632_), .B1(new_n643_), .B2(KEYINPUT69), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(KEYINPUT36), .A3(new_n631_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT69), .ZN(new_n646_));
  INV_X1    g445(.A(new_n632_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n639_), .A2(new_n646_), .A3(new_n647_), .A4(new_n642_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT70), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT70), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n644_), .A2(new_n645_), .A3(new_n651_), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT37), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(KEYINPUT37), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n628_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n283_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT38), .Z(new_n661_));
  INV_X1    g460(.A(new_n649_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n628_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n283_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT104), .Z(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(G1324gat));
  OAI21_X1  g465(.A(G8gat), .B1(new_n663_), .B2(new_n429_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(KEYINPUT39), .A3(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n659_), .A2(G8gat), .A3(new_n429_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n663_), .B2(new_n466_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n659_), .A2(G15gat), .A3(new_n466_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n663_), .B2(new_n462_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n659_), .A2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n462_), .B2(new_n684_), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n503_), .A2(new_n662_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n609_), .A2(new_n627_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n283_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n499_), .A2(new_n497_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n500_), .B1(new_n485_), .B2(new_n462_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT101), .B(new_n461_), .C1(new_n479_), .C2(new_n484_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n465_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n693_), .B(new_n657_), .C1(new_n698_), .C2(new_n464_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n503_), .B2(new_n658_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n502_), .A2(new_n466_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n464_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n705_), .A2(KEYINPUT107), .A3(new_n693_), .A4(new_n657_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n702_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n687_), .B(KEYINPUT106), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(KEYINPUT44), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n708_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n707_), .C2(new_n708_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n691_), .B(new_n709_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n692_), .B1(new_n716_), .B2(G29gat), .ZN(G1328gat));
  XNOR2_X1  g516(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n709_), .A2(new_n428_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n689_), .A2(G36gat), .A3(new_n429_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT45), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n721_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n718_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n726_), .B(new_n723_), .C1(new_n720_), .C2(G36gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1329gat));
  NOR2_X1   g527(.A1(new_n466_), .A2(new_n572_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n709_), .B(new_n729_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n572_), .B1(new_n689_), .B2(new_n466_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n690_), .B2(new_n461_), .ZN(new_n735_));
  OAI211_X1 g534(.A(G50gat), .B(new_n709_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(new_n461_), .ZN(G1331gat));
  INV_X1    g537(.A(new_n608_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n627_), .A2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n705_), .A2(new_n570_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n658_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n691_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n743_), .B2(new_n742_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(G57gat), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n741_), .A2(new_n662_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n283_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n746_), .B1(G57gat), .B2(new_n751_), .ZN(G1332gat));
  OR3_X1    g551(.A1(new_n742_), .A2(G64gat), .A3(new_n429_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n428_), .A3(new_n749_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G64gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G64gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1333gat));
  OR3_X1    g557(.A1(new_n742_), .A2(G71gat), .A3(new_n466_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n748_), .A2(new_n465_), .A3(new_n749_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G71gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n750_), .B2(new_n462_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT114), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n768_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n742_), .A2(G78gat), .A3(new_n462_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(G1335gat));
  INV_X1    g571(.A(new_n627_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n773_), .A2(new_n569_), .A3(new_n739_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n707_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(G85gat), .A3(new_n691_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n686_), .A2(new_n774_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n535_), .B1(new_n777_), .B2(new_n283_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n775_), .A2(G92gat), .A3(new_n428_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n536_), .B1(new_n777_), .B2(new_n429_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1337gat));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n707_), .A2(new_n465_), .A3(new_n774_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G99gat), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n466_), .A2(new_n532_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n777_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n783_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT51), .A3(new_n788_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n707_), .A2(new_n461_), .A3(new_n774_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G106gat), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n777_), .A2(G106gat), .A3(new_n462_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT116), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n465_), .A2(new_n691_), .A3(new_n462_), .A4(new_n429_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT120), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n607_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n598_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n566_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n553_), .A2(new_n554_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n555_), .A2(KEYINPUT55), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n553_), .A2(new_n812_), .A3(new_n554_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n563_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT55), .B(new_n557_), .C1(new_n546_), .C2(new_n552_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n817_), .A2(new_n818_), .B1(new_n554_), .B2(new_n553_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n563_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n809_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n605_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n599_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n592_), .A2(new_n593_), .ZN(new_n825_));
  MUX2_X1   g624(.A(new_n589_), .B(new_n825_), .S(new_n590_), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(new_n823_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n649_), .B1(new_n822_), .B2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n830_), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n565_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n815_), .B1(new_n814_), .B2(new_n563_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n820_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n829_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n662_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n832_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n831_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n565_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n827_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n566_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n828_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n846_), .A3(new_n657_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n662_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n822_), .A2(new_n829_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n851_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n662_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n847_), .A2(new_n850_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n841_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n850_), .A2(new_n852_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n830_), .B2(KEYINPUT57), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n838_), .A2(new_n832_), .A3(new_n839_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n855_), .A2(new_n858_), .A3(new_n859_), .A4(new_n847_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n854_), .A2(new_n627_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n740_), .A2(new_n569_), .A3(new_n658_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT54), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n806_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n830_), .A2(KEYINPUT57), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n627_), .B1(new_n853_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n805_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n245_), .A3(new_n608_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G113gat), .B1(new_n864_), .B2(new_n739_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1340gat));
  OAI211_X1 g674(.A(new_n570_), .B(new_n871_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G120gat), .ZN(new_n877_));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n864_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n878_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n877_), .A2(new_n880_), .A3(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1341gat));
  AOI21_X1  g684(.A(G127gat), .B1(new_n864_), .B2(new_n773_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT123), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n866_), .A2(G127gat), .A3(new_n773_), .A4(new_n871_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n872_), .A2(new_n890_), .A3(new_n658_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G134gat), .B1(new_n864_), .B2(new_n649_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  AOI21_X1  g692(.A(new_n428_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n466_), .A2(new_n461_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n283_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n608_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n226_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n569_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n227_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n627_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  NOR2_X1   g703(.A1(new_n897_), .A2(new_n662_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(G162gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n897_), .A2(new_n658_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(G162gat), .B2(new_n907_), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n350_), .A2(new_n461_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n869_), .A2(new_n428_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n289_), .B1(new_n911_), .B2(new_n739_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n912_), .A2(KEYINPUT62), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(new_n739_), .C1(new_n361_), .C2(new_n358_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(KEYINPUT62), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n861_), .A2(new_n863_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n917_), .A2(new_n428_), .A3(new_n909_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(G176gat), .A3(new_n570_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n290_), .B1(new_n910_), .B2(new_n569_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n918_), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n570_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(G1349gat));
  AOI21_X1  g723(.A(G183gat), .B1(new_n918_), .B2(new_n773_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n910_), .A2(new_n627_), .A3(new_n297_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n910_), .B2(new_n658_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n649_), .A2(new_n300_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n910_), .B2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n895_), .A2(new_n691_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n917_), .A2(new_n428_), .A3(new_n933_), .A4(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n608_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n376_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n569_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n374_), .ZN(G1353gat));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  AOI211_X1 g740(.A(new_n429_), .B(new_n934_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n942_), .A2(new_n773_), .A3(new_n933_), .A4(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n941_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n936_), .A2(new_n627_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n949_), .A2(KEYINPUT126), .A3(new_n944_), .A4(new_n946_), .ZN(new_n950_));
  OAI21_X1  g749(.A(KEYINPUT127), .B1(new_n949_), .B2(new_n944_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n952_), .B(new_n943_), .C1(new_n936_), .C2(new_n627_), .ZN(new_n953_));
  AOI22_X1  g752(.A1(new_n948_), .A2(new_n950_), .B1(new_n951_), .B2(new_n953_), .ZN(G1354gat));
  NOR2_X1   g753(.A1(new_n936_), .A2(new_n662_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(G218gat), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n936_), .A2(new_n658_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(G218gat), .B2(new_n957_), .ZN(G1355gat));
endmodule


