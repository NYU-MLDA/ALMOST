//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(KEYINPUT11), .B2(new_n202_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n205_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G231gat), .ZN(new_n217_));
  INV_X1    g016(.A(G233gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n216_), .B(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G127gat), .B(G155gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G183gat), .B(G211gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n225_), .B(KEYINPUT17), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n220_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n220_), .A2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n229_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n228_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G190gat), .B(G218gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G134gat), .B(G162gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT36), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT7), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n242_), .A2(new_n252_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G85gat), .ZN(new_n255_));
  INV_X1    g054(.A(G92gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G85gat), .A2(G92gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT65), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(KEYINPUT8), .A3(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n244_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n257_), .A2(KEYINPUT9), .A3(new_n258_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n258_), .A2(KEYINPUT9), .ZN(new_n269_));
  AND4_X1   g068(.A1(new_n251_), .A2(new_n267_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n262_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT8), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n264_), .A2(KEYINPUT66), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT66), .B1(new_n264_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G29gat), .B(G36gat), .Z(new_n277_));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT34), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT35), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(KEYINPUT35), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n264_), .A2(new_n273_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n279_), .B(KEYINPUT15), .ZN(new_n289_));
  AOI211_X1 g088(.A(new_n286_), .B(new_n287_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n280_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n280_), .B2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n241_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n240_), .B(KEYINPUT36), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT71), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n291_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT37), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT37), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n294_), .B(new_n298_), .C1(new_n300_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n237_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n276_), .A2(new_n208_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n276_), .A2(new_n208_), .ZN(new_n309_));
  OAI211_X1 g108(.A(G230gat), .B(G233gat), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n208_), .A2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n276_), .A2(new_n208_), .B1(new_n288_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n276_), .B2(new_n208_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G230gat), .A2(G233gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G120gat), .B(G148gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n310_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT13), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n324_), .B(new_n325_), .C1(KEYINPUT69), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n307_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT76), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT24), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n335_), .A2(new_n336_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G190gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT79), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT23), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT80), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT23), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n350_), .B1(new_n354_), .B2(KEYINPUT81), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n356_), .B(KEYINPUT23), .C1(new_n351_), .C2(new_n353_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n343_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n353_), .A3(KEYINPUT23), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n345_), .A2(new_n347_), .A3(G183gat), .A4(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n369_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G15gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT30), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n376_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(KEYINPUT84), .A3(new_n378_), .ZN(new_n382_));
  INV_X1    g181(.A(G120gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G113gat), .ZN(new_n384_));
  INV_X1    g183(.A(G113gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G120gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G134gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G127gat), .ZN(new_n391_));
  INV_X1    g190(.A(G127gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G134gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G113gat), .B(G120gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n389_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n389_), .B2(new_n396_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n381_), .A2(new_n382_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n382_), .A2(new_n401_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT2), .ZN(new_n406_));
  INV_X1    g205(.A(G141gat), .ZN(new_n407_));
  INV_X1    g206(.A(G148gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT85), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n415_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G141gat), .B(G148gat), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(KEYINPUT1), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n419_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n415_), .A2(KEYINPUT1), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n423_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n422_), .B(new_n427_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n428_));
  AND4_X1   g227(.A1(new_n409_), .A2(new_n412_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n421_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n389_), .A2(new_n396_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n397_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n389_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n436_), .A3(KEYINPUT4), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n431_), .A2(new_n434_), .A3(new_n438_), .A4(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT94), .Z(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n428_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G85gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT0), .B(G57gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n428_), .A2(new_n436_), .A3(KEYINPUT4), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n439_), .A2(new_n441_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n443_), .B(new_n448_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT27), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT19), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT21), .ZN(new_n459_));
  AND2_X1   g258(.A1(G197gat), .A2(G204gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G197gat), .A2(G204gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G197gat), .ZN(new_n463_));
  INV_X1    g262(.A(G204gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G197gat), .A2(G204gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT21), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G211gat), .B(G218gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n462_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n462_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT90), .B1(new_n467_), .B2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n362_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n366_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n340_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n342_), .B(KEYINPUT91), .Z(new_n479_));
  INV_X1    g278(.A(new_n341_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n473_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n358_), .A2(new_n473_), .A3(new_n368_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT20), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n458_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G8gat), .B(G36gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n492_));
  INV_X1    g291(.A(new_n473_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n369_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n458_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n477_), .A2(new_n473_), .A3(new_n481_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n485_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n491_), .B1(new_n485_), .B2(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n456_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n482_), .A2(new_n484_), .A3(new_n458_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n490_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT27), .A3(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n473_), .B1(KEYINPUT29), .B2(new_n431_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n510_), .B(new_n470_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n511_));
  INV_X1    g310(.A(G78gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G228gat), .A2(G233gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT89), .Z(new_n514_));
  AND3_X1   g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n244_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G78gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n520_));
  AOI21_X1  g319(.A(G106gat), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n244_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(G106gat), .A3(new_n520_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n508_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n523_), .A3(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G22gat), .B(G50gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n431_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT28), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT86), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n525_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT87), .B1(new_n536_), .B2(new_n509_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n528_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n526_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n455_), .B(new_n507_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT96), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n491_), .A2(KEYINPUT32), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n485_), .A2(new_n497_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n453_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n448_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n482_), .A2(new_n484_), .A3(new_n458_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n503_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT32), .B(new_n491_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n454_), .A2(KEYINPUT96), .A3(new_n554_), .A4(new_n546_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT95), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n442_), .A2(new_n443_), .A3(new_n448_), .A4(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n437_), .A2(new_n440_), .A3(new_n439_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n428_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n449_), .A3(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n485_), .A2(new_n497_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n490_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n453_), .A2(KEYINPUT95), .A3(new_n556_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n562_), .A2(new_n498_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n553_), .A2(new_n555_), .A3(new_n566_), .ZN(new_n567_));
  AND4_X1   g366(.A1(new_n523_), .A2(new_n522_), .A3(new_n538_), .A4(new_n526_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n538_), .B1(new_n537_), .B2(new_n526_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n534_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n540_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n405_), .B1(new_n543_), .B2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n541_), .A2(new_n542_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n402_), .A2(new_n455_), .A3(new_n403_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(new_n507_), .A3(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n279_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n215_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT77), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n289_), .A2(new_n215_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n577_), .A2(new_n215_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT78), .ZN(new_n589_));
  XOR2_X1   g388(.A(G169gat), .B(G197gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n576_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n333_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT97), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n454_), .A2(KEYINPUT98), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n454_), .A2(KEYINPUT98), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n210_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n299_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n237_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n576_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n592_), .A4(new_n331_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n455_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(G1324gat));
  NAND3_X1  g408(.A1(new_n596_), .A2(new_n211_), .A3(new_n506_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G8gat), .B1(new_n607_), .B2(new_n507_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT39), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n607_), .B2(new_n404_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT41), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n405_), .A2(new_n374_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n595_), .B2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n607_), .B2(new_n573_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n573_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n595_), .B2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n236_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n233_), .A2(new_n234_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n624_), .A2(new_n625_), .B1(new_n227_), .B2(new_n220_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n331_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n299_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n594_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n454_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n454_), .B(new_n506_), .C1(new_n570_), .C2(new_n540_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n567_), .A2(new_n540_), .A3(new_n570_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n404_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n573_), .A2(new_n507_), .A3(new_n574_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n305_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n632_), .B(KEYINPUT43), .C1(new_n637_), .C2(KEYINPUT101), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  NOR4_X1   g439(.A1(new_n626_), .A2(new_n627_), .A3(new_n593_), .A4(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n637_), .B2(new_n632_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n306_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n638_), .B(new_n641_), .C1(new_n643_), .C2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT104), .B1(new_n639_), .B2(KEYINPUT103), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n632_), .B1(new_n637_), .B2(KEYINPUT101), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT43), .B1(new_n644_), .B2(KEYINPUT102), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n648_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(new_n638_), .A3(new_n641_), .A4(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n599_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n631_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n630_), .A2(new_n658_), .A3(new_n506_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT45), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n655_), .A2(new_n506_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT105), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n507_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n658_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n662_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n662_), .A2(new_n665_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT106), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n662_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(KEYINPUT107), .A3(new_n670_), .A4(new_n660_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n673_), .A2(new_n678_), .ZN(G1329gat));
  XNOR2_X1  g478(.A(KEYINPUT109), .B(G43gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n629_), .B2(new_n404_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n655_), .A2(G43gat), .A3(new_n405_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n683_), .B2(new_n682_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g485(.A(new_n573_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G50gat), .B1(new_n630_), .B2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n655_), .B2(new_n689_), .ZN(G1331gat));
  NOR3_X1   g489(.A1(new_n576_), .A2(new_n592_), .A3(new_n331_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n605_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n455_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n307_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n599_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(G57gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n694_), .B2(new_n696_), .ZN(G1332gat));
  OAI21_X1  g496(.A(G64gat), .B1(new_n692_), .B2(new_n507_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT48), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n507_), .A2(G64gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n694_), .B2(new_n700_), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n692_), .B2(new_n404_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n404_), .A2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n694_), .B2(new_n704_), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n692_), .B2(new_n573_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n687_), .A2(new_n512_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n694_), .B2(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT110), .Z(G1335gat));
  NOR3_X1   g509(.A1(new_n626_), .A2(new_n592_), .A3(new_n331_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n652_), .A2(new_n638_), .A3(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT111), .Z(new_n713_));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n455_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n626_), .A2(new_n299_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n691_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n255_), .A3(new_n599_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1336gat));
  OAI21_X1  g518(.A(G92gat), .B1(new_n713_), .B2(new_n507_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n256_), .A3(new_n506_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1337gat));
  OAI21_X1  g521(.A(G99gat), .B1(new_n712_), .B2(new_n404_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n405_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n716_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT51), .ZN(G1338gat));
  OR2_X1    g525(.A1(new_n712_), .A2(new_n573_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(G106gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(KEYINPUT52), .A3(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n716_), .A2(G106gat), .A3(new_n573_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1339gat));
  AND2_X1   g538(.A1(new_n592_), .A2(new_n325_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n316_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n313_), .A2(new_n314_), .A3(KEYINPUT55), .A4(new_n315_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n323_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n747_), .B(new_n322_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT114), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n740_), .B(new_n751_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n587_), .A2(new_n591_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n584_), .A2(new_n585_), .A3(new_n580_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n578_), .A2(new_n579_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n591_), .A3(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n326_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n750_), .A2(new_n752_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT57), .B1(new_n759_), .B2(new_n299_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n757_), .A2(new_n325_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n761_), .B(KEYINPUT58), .C1(new_n746_), .C2(new_n748_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n306_), .A3(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n760_), .A2(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n759_), .A2(KEYINPUT57), .A3(new_n299_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n626_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n307_), .A2(new_n593_), .A3(new_n331_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT54), .Z(new_n772_));
  NOR2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n687_), .A2(new_n506_), .A3(new_n404_), .A4(new_n695_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G113gat), .B1(new_n776_), .B2(new_n592_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT115), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT118), .B1(new_n760_), .B2(new_n766_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n764_), .A2(new_n306_), .A3(new_n765_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n758_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n749_), .B2(KEYINPUT114), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n604_), .B1(new_n784_), .B2(new_n752_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n781_), .B(new_n782_), .C1(new_n785_), .C2(KEYINPUT57), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n780_), .A2(new_n769_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n772_), .B1(new_n787_), .B2(new_n237_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n779_), .B1(new_n788_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n782_), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n768_), .B1(new_n796_), .B2(KEYINPUT118), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n626_), .B1(new_n797_), .B2(new_n786_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT119), .B(new_n793_), .C1(new_n798_), .C2(new_n772_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n773_), .B2(new_n775_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n592_), .A2(G113gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT120), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n778_), .B1(new_n802_), .B2(new_n804_), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n801_), .B2(new_n331_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n383_), .B1(new_n331_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n776_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n383_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1341gat));
  OAI21_X1  g608(.A(G127gat), .B1(new_n801_), .B2(new_n237_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n776_), .A2(new_n392_), .A3(new_n626_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1342gat));
  OAI21_X1  g611(.A(G134gat), .B1(new_n801_), .B2(new_n305_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n776_), .A2(new_n390_), .A3(new_n604_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT121), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n817_), .A3(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1343gat));
  NAND3_X1  g618(.A1(new_n404_), .A2(new_n507_), .A3(new_n599_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n773_), .A2(new_n573_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n592_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n627_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n626_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  AOI21_X1  g627(.A(G162gat), .B1(new_n821_), .B2(new_n604_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n306_), .A2(G162gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT122), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n821_), .B2(new_n831_), .ZN(G1347gat));
  NOR4_X1   g631(.A1(new_n687_), .A2(new_n507_), .A3(new_n404_), .A4(new_n599_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n592_), .B(new_n833_), .C1(new_n798_), .C2(new_n772_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n835_), .A3(G169gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n834_), .B2(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n833_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n788_), .A2(new_n593_), .A3(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT123), .B(new_n838_), .C1(new_n841_), .C2(new_n335_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT22), .B(G169gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT124), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n837_), .A2(new_n838_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n837_), .A2(new_n838_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n847_), .B(new_n848_), .C1(new_n849_), .C2(new_n836_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(G1348gat));
  NOR2_X1   g650(.A1(new_n773_), .A2(new_n840_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(G176gat), .A3(new_n627_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n788_), .A2(new_n331_), .A3(new_n840_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(G176gat), .B2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT125), .ZN(G1349gat));
  AOI21_X1  g655(.A(G183gat), .B1(new_n852_), .B2(new_n626_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n788_), .A2(new_n840_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n626_), .A2(new_n479_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT126), .ZN(G1350gat));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n341_), .A3(new_n604_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n788_), .A2(new_n305_), .A3(new_n840_), .ZN(new_n863_));
  INV_X1    g662(.A(G190gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1351gat));
  NAND4_X1  g664(.A1(new_n687_), .A2(new_n455_), .A3(new_n506_), .A4(new_n404_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n773_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n592_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n627_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g670(.A(new_n237_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT127), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n875_));
  INV_X1    g674(.A(G211gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n874_), .B(new_n877_), .ZN(G1354gat));
  INV_X1    g677(.A(new_n867_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G218gat), .B1(new_n879_), .B2(new_n305_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n299_), .A2(G218gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n879_), .B2(new_n881_), .ZN(G1355gat));
endmodule


