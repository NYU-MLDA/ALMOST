//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT13), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(KEYINPUT13), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G120gat), .B(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT5), .B(G176gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n209_), .B(new_n210_), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G71gat), .B(G78gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n215_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(KEYINPUT11), .C2(new_n213_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(KEYINPUT11), .A3(new_n219_), .A4(new_n213_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT67), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240_));
  INV_X1    g039(.A(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n236_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n231_), .A2(new_n235_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n237_), .B2(new_n238_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n241_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(KEYINPUT65), .A3(new_n232_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n230_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n256_));
  OAI22_X1  g055(.A1(new_n243_), .A2(new_n244_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(new_n255_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n241_), .A2(new_n236_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT9), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT10), .B(G99gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT64), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n258_), .B(new_n261_), .C1(new_n263_), .C2(G106gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n224_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n224_), .A2(new_n265_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n258_), .A2(new_n231_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n245_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n254_), .A2(new_n232_), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n247_), .A2(new_n248_), .B1(new_n272_), .B2(new_n230_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n270_), .A2(new_n271_), .B1(new_n273_), .B2(KEYINPUT8), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT10), .B(G99gat), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT64), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n262_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(G106gat), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n258_), .A2(new_n261_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT70), .B1(new_n274_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n257_), .A2(new_n283_), .A3(new_n264_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT12), .A3(new_n224_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G230gat), .A2(G233gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n269_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n267_), .B1(new_n290_), .B2(new_n266_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n266_), .A2(new_n290_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n212_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n266_), .A2(new_n290_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n224_), .B2(new_n265_), .ZN(new_n297_));
  OAI211_X1 g096(.A(G230gat), .B(G233gat), .C1(new_n297_), .C2(new_n292_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n288_), .A3(new_n211_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n299_), .A3(KEYINPUT71), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT71), .B1(new_n295_), .B2(new_n299_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n205_), .B(new_n206_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(new_n299_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT13), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(KEYINPUT72), .A3(new_n307_), .A4(new_n300_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G169gat), .B(G197gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G141gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G229gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT77), .B(G8gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT14), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G1gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(KEYINPUT14), .A2(G1gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G8gat), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n318_), .A2(G1gat), .B1(new_n315_), .B2(new_n320_), .ZN(new_n324_));
  INV_X1    g123(.A(G8gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G29gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G43gat), .B(G50gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n314_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n322_), .A2(G8gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n324_), .A2(new_n325_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n329_), .B(KEYINPUT15), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n331_), .B(new_n313_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n312_), .B1(new_n341_), .B2(KEYINPUT79), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(KEYINPUT79), .B2(new_n341_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT80), .B1(new_n340_), .B2(new_n312_), .ZN(new_n344_));
  AND4_X1   g143(.A1(KEYINPUT80), .A2(new_n334_), .A3(new_n339_), .A4(new_n312_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G231gat), .A2(G233gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n337_), .B(new_n348_), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(new_n224_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n351_));
  XNOR2_X1  g150(.A(G127gat), .B(G155gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G183gat), .B(G211gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n350_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n350_), .A2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G190gat), .B(G218gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G134gat), .B(G162gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT36), .ZN(new_n365_));
  INV_X1    g164(.A(new_n338_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n285_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G232gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT74), .B1(new_n370_), .B2(KEYINPUT35), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n370_), .A2(KEYINPUT35), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(KEYINPUT74), .A3(KEYINPUT35), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n265_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n330_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n367_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n338_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n374_), .B(new_n373_), .C1(new_n265_), .C2(new_n329_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n371_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n364_), .A2(KEYINPUT36), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n378_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n365_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n360_), .A2(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n309_), .A2(new_n347_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT30), .B(G15gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(KEYINPUT31), .Z(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401_));
  INV_X1    g200(.A(G183gat), .ZN(new_n402_));
  INV_X1    g201(.A(G190gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT24), .ZN(new_n405_));
  INV_X1    g204(.A(G169gat), .ZN(new_n406_));
  INV_X1    g205(.A(G176gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n404_), .A2(new_n408_), .A3(KEYINPUT83), .A4(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n407_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT26), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(KEYINPUT82), .B(KEYINPUT26), .C1(new_n418_), .C2(new_n419_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n403_), .A2(KEYINPUT26), .ZN(new_n424_));
  OR2_X1    g223(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n414_), .A2(new_n417_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT22), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(G169gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(G176gat), .B1(new_n431_), .B2(G169gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n406_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n416_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT85), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n438_), .A3(new_n416_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n402_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n429_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G71gat), .B(G99gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G43gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n400_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n400_), .A2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451_));
  INV_X1    g250(.A(G92gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT18), .B(G64gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT19), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n208_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(G197gat), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G197gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n208_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n461_), .A2(new_n465_), .A3(KEYINPUT21), .A4(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(G197gat), .B1(new_n463_), .B2(new_n464_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT21), .B1(new_n466_), .B2(new_n208_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n460_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT21), .B1(new_n465_), .B2(new_n467_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n468_), .B(KEYINPUT93), .C1(new_n471_), .C2(new_n472_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n429_), .A4(new_n442_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT20), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT22), .B(G169gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n407_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n416_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT95), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n402_), .A2(new_n403_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n404_), .A2(new_n409_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n489_), .A3(new_n416_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n483_), .A2(new_n487_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT26), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n427_), .B1(new_n492_), .B2(G190gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n410_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n417_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n478_), .A2(new_n479_), .B1(new_n473_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n477_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n459_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT20), .B1(new_n496_), .B2(new_n473_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n475_), .A2(new_n476_), .B1(new_n429_), .B2(new_n442_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n458_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n456_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n477_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT94), .B1(new_n477_), .B2(KEYINPUT20), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n473_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n504_), .B(new_n455_), .C1(new_n509_), .C2(new_n459_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT27), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n478_), .A2(new_n479_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n498_), .A3(new_n507_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n502_), .B1(new_n514_), .B2(new_n458_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n515_), .B2(new_n455_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n513_), .A2(new_n498_), .A3(new_n459_), .A4(new_n507_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n458_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n455_), .B(KEYINPUT98), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n511_), .A2(new_n512_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n523_));
  INV_X1    g322(.A(G141gat), .ZN(new_n524_));
  INV_X1    g323(.A(G148gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G155gat), .A2(G162gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT1), .Z(new_n531_));
  NOR2_X1   g330(.A1(G155gat), .A2(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT88), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT2), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT3), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT3), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(G141gat), .B2(G148gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n539_), .A2(new_n540_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT90), .A3(new_n536_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n533_), .A2(new_n530_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n534_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n523_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n552_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n557_));
  NOR4_X1   g356(.A1(new_n557_), .A2(KEYINPUT28), .A3(new_n534_), .A4(KEYINPUT29), .ZN(new_n558_));
  OAI21_X1  g357(.A(G22gat), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT90), .B1(new_n549_), .B2(new_n536_), .ZN(new_n560_));
  AND4_X1   g359(.A1(KEYINPUT90), .A2(new_n536_), .A3(new_n541_), .A4(new_n545_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n553_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n534_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT28), .B1(new_n564_), .B2(KEYINPUT29), .ZN(new_n565_));
  INV_X1    g364(.A(G22gat), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n554_), .A2(new_n523_), .A3(new_n555_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G50gat), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n559_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n559_), .B2(new_n568_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n475_), .A2(new_n476_), .B1(G228gat), .B2(G233gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT29), .B1(new_n557_), .B2(new_n534_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G228gat), .A2(G233gat), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n575_), .B2(new_n473_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G78gat), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G78gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n575_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n473_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n564_), .B2(KEYINPUT29), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n580_), .B(new_n581_), .C1(new_n583_), .C2(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n227_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(G106gat), .A3(new_n584_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n572_), .A2(new_n573_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n559_), .A2(new_n568_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G50gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n559_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n573_), .ZN(new_n593_));
  AOI21_X1  g392(.A(G106gat), .B1(new_n579_), .B2(new_n584_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n394_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n395_), .B1(new_n557_), .B2(new_n534_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(KEYINPUT4), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT4), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n564_), .A2(new_n603_), .A3(new_n395_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G225gat), .A2(G233gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G1gat), .B(G29gat), .ZN(new_n609_));
  INV_X1    g408(.A(G85gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT0), .B(G57gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  AOI21_X1  g412(.A(new_n607_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617_));
  INV_X1    g416(.A(new_n613_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n606_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(new_n614_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT97), .B(new_n618_), .C1(new_n619_), .C2(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n522_), .A2(new_n596_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n455_), .A2(KEYINPUT32), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n625_), .B(new_n504_), .C1(new_n509_), .C2(new_n459_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n519_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n621_), .A2(new_n622_), .A3(new_n626_), .A4(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n620_), .A2(KEYINPUT33), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n631_), .B(new_n618_), .C1(new_n619_), .C2(new_n614_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n600_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n613_), .B(new_n634_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n633_), .A2(new_n635_), .A3(new_n510_), .A4(new_n503_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n596_), .B1(new_n629_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n450_), .B1(new_n624_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n521_), .A2(KEYINPUT27), .A3(new_n510_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT27), .B1(new_n503_), .B2(new_n510_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n515_), .A2(new_n455_), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n456_), .B(new_n502_), .C1(new_n514_), .C2(new_n458_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n512_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n516_), .A2(new_n521_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(KEYINPUT99), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n588_), .A2(new_n595_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n623_), .A2(new_n449_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n642_), .A2(new_n647_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n638_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n388_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n623_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n202_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n347_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT100), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT37), .B1(new_n385_), .B2(KEYINPUT75), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT76), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n372_), .B1(new_n367_), .B2(new_n377_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n379_), .A2(new_n380_), .A3(new_n371_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n382_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n378_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n664_), .B2(new_n365_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n365_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT76), .B(new_n666_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n658_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n386_), .A2(KEYINPUT76), .ZN(new_n669_));
  INV_X1    g468(.A(new_n658_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n659_), .A3(new_n365_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n360_), .B1(new_n668_), .B2(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n309_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n657_), .A2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(new_n202_), .A3(new_n654_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n655_), .B1(new_n676_), .B2(KEYINPUT38), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(KEYINPUT101), .A3(KEYINPUT38), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n202_), .A3(new_n654_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT38), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n677_), .B1(new_n678_), .B2(new_n682_), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n642_), .A2(new_n647_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n316_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n684_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n652_), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1325gat));
  INV_X1    g491(.A(G15gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n675_), .A2(new_n693_), .A3(new_n449_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n653_), .B2(new_n449_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n697_), .A3(new_n698_), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n596_), .A2(new_n566_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT103), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n675_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G22gat), .B1(new_n652_), .B2(new_n648_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n360_), .A2(new_n386_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n309_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n657_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n654_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n309_), .A2(new_n347_), .A3(new_n360_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n668_), .A2(new_n672_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n633_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n503_), .A2(new_n635_), .A3(new_n510_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n629_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n648_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n522_), .A2(new_n596_), .A3(new_n623_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n449_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AND4_X1   g518(.A1(new_n648_), .A2(new_n642_), .A3(new_n647_), .A4(new_n649_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n713_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n668_), .A2(KEYINPUT104), .A3(new_n672_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT43), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n723_), .B(new_n713_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n711_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT44), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n729_), .B1(new_n727_), .B2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n654_), .A2(G29gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n710_), .B1(new_n733_), .B2(new_n734_), .ZN(G1328gat));
  NOR2_X1   g534(.A1(new_n687_), .A2(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n657_), .A2(new_n708_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n657_), .A2(new_n739_), .A3(new_n708_), .A4(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n711_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n723_), .B1(new_n651_), .B2(new_n713_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n726_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n742_), .B(new_n732_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n745_), .B(new_n684_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT107), .B1(new_n746_), .B2(G36gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n741_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n741_), .B(KEYINPUT46), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1329gat));
  NAND3_X1  g552(.A1(new_n733_), .A2(G43gat), .A3(new_n449_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n657_), .A2(new_n449_), .A3(new_n708_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT108), .B(G43gat), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT47), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1330gat));
  NAND2_X1  g561(.A1(new_n596_), .A2(new_n569_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT109), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n709_), .A2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n733_), .A2(new_n596_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n569_), .ZN(G1331gat));
  INV_X1    g566(.A(G57gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n347_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n309_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n651_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n673_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n772_), .B2(new_n623_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n387_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n654_), .A2(G57gat), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n773_), .A2(KEYINPUT110), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(KEYINPUT110), .B2(new_n773_), .ZN(G1332gat));
  OR3_X1    g576(.A1(new_n772_), .A2(G64gat), .A3(new_n687_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n684_), .A3(new_n387_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(G64gat), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(G64gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  OR3_X1    g583(.A1(new_n772_), .A2(G71gat), .A3(new_n450_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n449_), .A3(new_n387_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(G71gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n786_), .B2(G71gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(G1334gat));
  NAND3_X1  g590(.A1(new_n771_), .A2(new_n596_), .A3(new_n387_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(G78gat), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n792_), .B2(G78gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n596_), .A2(new_n580_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n795_), .A2(new_n796_), .B1(new_n772_), .B2(new_n797_), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n771_), .A2(new_n707_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G85gat), .B1(new_n800_), .B2(new_n654_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n770_), .A2(new_n769_), .A3(new_n360_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n623_), .A2(new_n610_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(G1336gat));
  AOI21_X1  g604(.A(G92gat), .B1(new_n800_), .B2(new_n684_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n684_), .A2(G92gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT111), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n803_), .B2(new_n808_), .ZN(G1337gat));
  NAND2_X1  g608(.A1(new_n803_), .A2(new_n449_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n810_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT112), .B1(new_n810_), .B2(G99gat), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n450_), .A2(new_n263_), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n811_), .A2(new_n812_), .B1(new_n799_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n814_), .B(new_n816_), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n803_), .A2(new_n596_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(G106gat), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT52), .B(new_n227_), .C1(new_n803_), .C2(new_n596_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n596_), .A2(new_n227_), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n820_), .A2(new_n821_), .B1(new_n799_), .B2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g623(.A(new_n287_), .B1(new_n269_), .B2(new_n286_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n288_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n269_), .A2(new_n286_), .A3(KEYINPUT55), .A4(new_n287_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n211_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n289_), .A2(new_n294_), .A3(new_n212_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n833_), .A3(new_n347_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n329_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n314_), .B1(new_n835_), .B2(new_n331_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n836_), .A2(KEYINPUT114), .A3(new_n312_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n331_), .B(new_n314_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT114), .B1(new_n836_), .B2(new_n312_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT115), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n840_), .B(new_n843_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n300_), .A3(new_n306_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n386_), .B1(new_n834_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT57), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n831_), .A2(new_n845_), .A3(new_n833_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n831_), .A2(new_n845_), .A3(new_n833_), .A4(KEYINPUT58), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n713_), .A3(new_n852_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n854_));
  OAI211_X1 g653(.A(new_n848_), .B(new_n853_), .C1(new_n847_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n360_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n309_), .A2(new_n769_), .A3(new_n673_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT54), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n309_), .A2(new_n859_), .A3(new_n769_), .A4(new_n673_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n684_), .A2(new_n623_), .A3(new_n596_), .A4(new_n450_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n347_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n853_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n853_), .B(KEYINPUT117), .C1(new_n847_), .C2(new_n854_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n848_), .A3(new_n871_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n872_), .A2(new_n360_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n863_), .A2(new_n867_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n865_), .A2(new_n867_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n347_), .A2(G113gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n866_), .B1(new_n876_), .B2(new_n877_), .ZN(G1340gat));
  XOR2_X1   g677(.A(KEYINPUT118), .B(G120gat), .Z(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT60), .B1(new_n770_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n770_), .B1(new_n864_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n875_), .B2(new_n882_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n864_), .A2(new_n881_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(KEYINPUT60), .B2(new_n884_), .ZN(G1341gat));
  INV_X1    g684(.A(new_n360_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G127gat), .B1(new_n865_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(G127gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT119), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n876_), .B2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n865_), .B2(new_n386_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n713_), .A2(G134gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n876_), .B2(new_n892_), .ZN(G1343gat));
  AOI22_X1  g692(.A1(new_n855_), .A2(new_n360_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n687_), .A2(new_n654_), .A3(new_n450_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n648_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n347_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT120), .B(G141gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n770_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT121), .B(G148gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  NAND2_X1  g701(.A1(new_n896_), .A2(new_n886_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n896_), .B2(new_n386_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n713_), .A2(G162gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n896_), .B2(new_n907_), .ZN(G1347gat));
  NAND3_X1  g707(.A1(new_n684_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n873_), .A2(new_n769_), .A3(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n910_), .A2(new_n406_), .A3(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n910_), .B2(new_n406_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n873_), .A2(new_n909_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n347_), .A2(new_n480_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT123), .Z(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n913_), .A2(new_n914_), .A3(new_n918_), .ZN(G1348gat));
  NOR4_X1   g718(.A1(new_n894_), .A2(new_n407_), .A3(new_n309_), .A4(new_n909_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n915_), .A2(new_n770_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n407_), .ZN(G1349gat));
  OR3_X1    g721(.A1(new_n894_), .A2(new_n360_), .A3(new_n909_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(KEYINPUT124), .ZN(new_n924_));
  AOI21_X1  g723(.A(G183gat), .B1(new_n923_), .B2(KEYINPUT124), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n886_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n915_), .B2(new_n926_), .ZN(G1350gat));
  NOR2_X1   g726(.A1(new_n492_), .A2(G190gat), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n424_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n915_), .A2(new_n386_), .A3(new_n929_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n873_), .A2(new_n712_), .A3(new_n909_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n403_), .ZN(G1351gat));
  AOI21_X1  g731(.A(new_n648_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n684_), .A2(new_n623_), .A3(new_n450_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n933_), .B2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n894_), .A2(new_n937_), .A3(new_n648_), .A4(new_n934_), .ZN(new_n938_));
  OAI211_X1 g737(.A(G197gat), .B(new_n347_), .C1(new_n936_), .C2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n862_), .A2(new_n596_), .A3(new_n935_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n937_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n933_), .A2(KEYINPUT125), .A3(new_n935_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n945_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n347_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n347_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n466_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n941_), .A2(new_n946_), .A3(new_n948_), .ZN(G1352gat));
  AOI21_X1  g748(.A(new_n309_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n463_), .A2(new_n464_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n950_), .B2(new_n208_), .ZN(G1353gat));
  OR2_X1    g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n945_), .B2(new_n886_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n360_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n956_));
  XOR2_X1   g755(.A(KEYINPUT63), .B(G211gat), .Z(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(G1354gat));
  AOI21_X1  g757(.A(G218gat), .B1(new_n945_), .B2(new_n386_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n713_), .A2(G218gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT127), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n945_), .B2(new_n961_), .ZN(G1355gat));
endmodule


