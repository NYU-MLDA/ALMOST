//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_;
  INV_X1    g000(.A(G127gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(G120gat), .A3(new_n205_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT80), .B(G113gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT82), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n217_), .A2(KEYINPUT83), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(new_n219_), .A3(KEYINPUT1), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(G155gat), .A4(G162gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n227_), .B2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(KEYINPUT84), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT2), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(KEYINPUT84), .A3(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G155gat), .B(G162gat), .Z(new_n238_));
  AOI22_X1  g037(.A1(new_n224_), .A2(new_n229_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n213_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n211_), .A2(new_n212_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n224_), .A2(new_n229_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n245_), .A3(KEYINPUT4), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(KEYINPUT4), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n252_));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n240_), .A2(new_n245_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n249_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n258_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(G197gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT87), .B1(new_n273_), .B2(G204gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(G204gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n268_), .B(new_n272_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n267_), .B1(new_n280_), .B2(new_n268_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n277_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT25), .B(G183gat), .Z(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT26), .B(G190gat), .Z(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT24), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT77), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n289_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n284_), .B1(new_n287_), .B2(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n293_), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT77), .B1(new_n290_), .B2(new_n291_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT24), .B(new_n288_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(KEYINPUT91), .C1(new_n285_), .C2(new_n286_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT23), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n292_), .A2(KEYINPUT24), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT92), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT92), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n303_), .B(new_n307_), .C1(KEYINPUT24), .C2(new_n292_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n297_), .A2(new_n301_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n288_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n291_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT93), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  INV_X1    g113(.A(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n303_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n303_), .B2(new_n316_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n283_), .B1(new_n309_), .B2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT76), .B(G190gat), .Z(new_n321_));
  OAI21_X1  g120(.A(new_n303_), .B1(G183gat), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n312_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n294_), .A2(new_n295_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n300_), .B(new_n303_), .C1(KEYINPUT24), .C2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n326_));
  OR2_X1    g125(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n285_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT20), .B1(new_n329_), .B2(new_n282_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n266_), .B1(new_n320_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n309_), .A2(new_n283_), .A3(new_n319_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n266_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n282_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n332_), .A2(KEYINPUT20), .A3(new_n333_), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G64gat), .B(G92gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n331_), .A2(new_n341_), .A3(new_n335_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT27), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n320_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n330_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n333_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT99), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT99), .A4(new_n333_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n332_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT98), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n354_), .A2(new_n355_), .B1(new_n282_), .B2(new_n329_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n332_), .A2(KEYINPUT98), .A3(new_n353_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n333_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n342_), .B1(new_n352_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n344_), .A2(KEYINPUT27), .ZN(new_n360_));
  AOI211_X1 g159(.A(new_n264_), .B(new_n345_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT31), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n329_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n323_), .B(new_n363_), .C1(new_n325_), .C2(new_n328_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G71gat), .B(G99gat), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT78), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n213_), .A2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(new_n211_), .A2(new_n212_), .A3(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G15gat), .B(G43gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n380_), .A3(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n369_), .A2(new_n379_), .A3(new_n371_), .A4(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n239_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n239_), .B2(new_n389_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n388_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n283_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n282_), .A2(KEYINPUT88), .ZN(new_n401_));
  INV_X1    g200(.A(G228gat), .ZN(new_n402_));
  INV_X1    g201(.A(G233gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n403_), .A2(KEYINPUT86), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(KEYINPUT86), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n282_), .B1(new_n239_), .B2(new_n389_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G78gat), .B(G106gat), .Z(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n398_), .B(new_n412_), .C1(new_n413_), .C2(KEYINPUT89), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(KEYINPUT89), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT90), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n398_), .A2(new_n412_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n410_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n411_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n413_), .A2(KEYINPUT89), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n417_), .A2(new_n422_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n398_), .B1(new_n420_), .B2(new_n412_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n386_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n427_), .B(new_n385_), .C1(new_n416_), .C2(new_n425_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n361_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n343_), .A2(new_n344_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT95), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n343_), .A2(KEYINPUT95), .A3(new_n344_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n263_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT33), .B(new_n260_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n248_), .A2(new_n250_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n256_), .B1(new_n257_), .B2(new_n249_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n438_), .B(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n352_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n358_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n264_), .B1(new_n443_), .B2(new_n336_), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n436_), .A2(new_n442_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n426_), .A2(new_n428_), .A3(new_n385_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n431_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G1gat), .A2(G8gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT14), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n456_), .B(KEYINPUT71), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G29gat), .B(G36gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G43gat), .B(G50gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n470_), .A2(new_n473_), .A3(KEYINPUT74), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT74), .B1(new_n470_), .B2(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n470_), .A2(new_n473_), .A3(KEYINPUT15), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n470_), .B2(new_n473_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n464_), .B(new_n466_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT75), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n477_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n464_), .B(new_n466_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n477_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n455_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n455_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n452_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT100), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT100), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n452_), .A2(new_n496_), .A3(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT11), .ZN(new_n499_));
  INV_X1    g298(.A(G57gat), .ZN(new_n500_));
  INV_X1    g299(.A(G64gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G57gat), .A2(G64gat), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  AND2_X1   g306(.A1(G71gat), .A2(G78gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G71gat), .A2(G78gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n505_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(G57gat), .A2(G64gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G57gat), .A2(G64gat), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G71gat), .B(G78gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT65), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n504_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G231gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n403_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n467_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n467_), .A2(new_n523_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n521_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n526_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n511_), .A2(new_n512_), .A3(new_n505_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n504_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n531_), .A3(new_n524_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n527_), .A2(new_n532_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(KEYINPUT73), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n539_), .B(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n542_), .B2(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n534_), .A2(new_n544_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(G106gat), .ZN(new_n551_));
  INV_X1    g350(.A(G99gat), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(KEYINPUT10), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(KEYINPUT10), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT64), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n555_), .B(new_n560_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n552_), .A3(new_n551_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n558_), .A3(new_n559_), .A4(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT8), .ZN(new_n575_));
  INV_X1    g374(.A(new_n561_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n565_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n570_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT8), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n470_), .A2(new_n473_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n587_), .A3(new_n570_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT35), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(KEYINPUT35), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595_));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n581_), .A2(KEYINPUT35), .A3(new_n590_), .A4(new_n588_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n598_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n594_), .B2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT70), .B1(new_n602_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n594_), .A2(new_n600_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n601_), .B1(new_n609_), .B2(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n550_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n614_));
  OR2_X1    g413(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n271_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT5), .B(G176gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n580_), .B1(new_n520_), .B2(new_n513_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT67), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n585_), .B(new_n570_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT67), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n622_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT12), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n531_), .B(new_n580_), .C1(KEYINPUT66), .C2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n580_), .B2(KEYINPUT66), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n580_), .A2(new_n520_), .A3(new_n513_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n624_), .A2(new_n627_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n625_), .A2(new_n631_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n622_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n620_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n629_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n626_), .B1(new_n625_), .B2(new_n622_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n555_), .A2(new_n560_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n568_), .A2(new_n569_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n583_), .A2(new_n584_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT67), .B(new_n623_), .C1(new_n641_), .C2(new_n521_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n637_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n635_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n619_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n636_), .A2(new_n645_), .A3(KEYINPUT68), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT68), .B1(new_n636_), .B2(new_n645_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n614_), .B(new_n615_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n636_), .A2(new_n645_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT68), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n652_), .A2(KEYINPUT69), .A3(KEYINPUT13), .A4(new_n646_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n649_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n498_), .A2(new_n613_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n264_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(G1gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n653_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n613_), .A4(new_n657_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(KEYINPUT38), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n654_), .A2(new_n665_), .A3(new_n549_), .A4(new_n493_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n610_), .B1(new_n431_), .B2(new_n451_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n649_), .A2(new_n653_), .A3(new_n549_), .A4(new_n493_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT102), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n656_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n664_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT38), .B1(new_n659_), .B2(new_n663_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT103), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n659_), .A2(new_n663_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n671_), .A4(new_n664_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(G1324gat));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n359_), .A2(new_n360_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n345_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(G8gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n681_), .B1(new_n655_), .B2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n661_), .A2(KEYINPUT104), .A3(new_n613_), .A4(new_n686_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n666_), .A2(new_n667_), .A3(new_n684_), .A4(new_n669_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n691_), .B2(G8gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT39), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT106), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(G8gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n691_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(KEYINPUT106), .A3(new_n695_), .A4(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT39), .B1(new_n692_), .B2(new_n693_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n690_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT40), .B(new_n690_), .C1(new_n696_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1325gat));
  OR3_X1    g507(.A1(new_n655_), .A2(G15gat), .A3(new_n385_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G15gat), .B1(new_n670_), .B2(new_n385_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT41), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT41), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n711_), .A3(new_n712_), .ZN(G1326gat));
  NAND2_X1  g512(.A1(new_n426_), .A2(new_n428_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G22gat), .B1(new_n670_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT42), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(G22gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT107), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n655_), .B2(new_n719_), .ZN(G1327gat));
  NOR3_X1   g519(.A1(new_n660_), .A2(new_n549_), .A3(new_n492_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n452_), .A2(new_n612_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT43), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT43), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n721_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n264_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G29gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n610_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n549_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n661_), .A2(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n656_), .A2(G29gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1328gat));
  NOR2_X1   g534(.A1(new_n685_), .A2(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n661_), .A2(new_n732_), .A3(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT45), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n684_), .A3(new_n728_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n740_), .A3(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  NAND3_X1  g544(.A1(new_n727_), .A2(new_n386_), .A3(new_n728_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G43gat), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n733_), .A2(G43gat), .A3(new_n385_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(KEYINPUT47), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1330gat));
  NAND3_X1  g552(.A1(new_n727_), .A2(new_n714_), .A3(new_n728_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G50gat), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n715_), .A2(G50gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n733_), .B2(new_n756_), .ZN(G1331gat));
  AOI21_X1  g556(.A(new_n493_), .B1(new_n431_), .B2(new_n451_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n660_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n550_), .A2(new_n610_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(G57gat), .A3(new_n264_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n660_), .A2(new_n613_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT108), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT108), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n758_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n264_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n500_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(KEYINPUT109), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n763_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n501_), .B1(new_n761_), .B2(new_n684_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT48), .Z(new_n775_));
  NAND3_X1  g574(.A1(new_n767_), .A2(new_n501_), .A3(new_n684_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1333gat));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n767_), .A2(new_n778_), .A3(new_n386_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n761_), .A2(new_n386_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(G71gat), .ZN(new_n782_));
  AOI211_X1 g581(.A(KEYINPUT49), .B(new_n778_), .C1(new_n761_), .C2(new_n386_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT111), .ZN(G1334gat));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n761_), .B2(new_n714_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT50), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n767_), .A2(new_n786_), .A3(new_n714_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1335gat));
  NAND3_X1  g589(.A1(new_n759_), .A2(KEYINPUT112), .A3(new_n732_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n758_), .A2(new_n660_), .A3(new_n732_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n264_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n723_), .A2(new_n724_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n654_), .A2(new_n549_), .A3(new_n493_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n264_), .A2(G85gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(G1336gat));
  AOI21_X1  g600(.A(G92gat), .B1(new_n795_), .B2(new_n684_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n684_), .A2(G92gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n799_), .B2(new_n803_), .ZN(G1337gat));
  OAI211_X1 g603(.A(new_n386_), .B(new_n798_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(G99gat), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n805_), .B2(G99gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT115), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n553_), .A2(new_n554_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n385_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT51), .B1(new_n810_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n809_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n807_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n814_), .B(KEYINPUT114), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(KEYINPUT115), .A4(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(G1338gat));
  NAND3_X1  g622(.A1(new_n795_), .A2(new_n551_), .A3(new_n714_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n714_), .B(new_n798_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(new_n826_), .A3(G106gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n825_), .B2(G106gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT53), .ZN(G1339gat));
  AND4_X1   g629(.A1(new_n549_), .A2(new_n611_), .A3(new_n608_), .A4(new_n492_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n653_), .A3(new_n649_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n477_), .A2(new_n480_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n477_), .A2(new_n837_), .A3(new_n480_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n482_), .A3(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n477_), .A2(new_n486_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n839_), .B(new_n455_), .C1(new_n840_), .C2(new_n482_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n491_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n652_), .B2(new_n646_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n642_), .A2(new_n638_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n632_), .A2(new_n629_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n637_), .B(KEYINPUT55), .C1(new_n638_), .C2(new_n642_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n623_), .B1(new_n847_), .B2(new_n621_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n851_), .B2(new_n620_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(KEYINPUT116), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n851_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n620_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n633_), .A2(new_n635_), .A3(new_n620_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n492_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n844_), .B1(new_n854_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n731_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n621_), .B1(new_n632_), .B2(new_n629_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n633_), .A2(KEYINPUT55), .B1(new_n622_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n849_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n620_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n620_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n855_), .A2(new_n857_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n843_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n860_), .B1(new_n873_), .B2(new_n610_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n612_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n842_), .A2(new_n856_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n876_), .B(KEYINPUT58), .C1(new_n852_), .C2(new_n853_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n862_), .A2(new_n874_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n834_), .B1(new_n882_), .B2(new_n550_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n430_), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n883_), .A2(new_n656_), .A3(new_n884_), .A4(new_n684_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G113gat), .B1(new_n885_), .B2(new_n493_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n883_), .A2(new_n656_), .A3(new_n684_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n430_), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n885_), .A2(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n493_), .A2(G113gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n886_), .B1(new_n894_), .B2(new_n895_), .ZN(G1340gat));
  OAI21_X1  g695(.A(new_n207_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n885_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n207_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n654_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n207_), .ZN(G1341gat));
  AOI21_X1  g699(.A(G127gat), .B1(new_n885_), .B2(new_n549_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n550_), .A2(new_n202_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n894_), .B2(new_n902_), .ZN(G1342gat));
  AOI21_X1  g702(.A(G134gat), .B1(new_n885_), .B2(new_n610_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n875_), .A2(new_n203_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n894_), .B2(new_n905_), .ZN(G1343gat));
  AND2_X1   g705(.A1(new_n887_), .A2(new_n429_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n493_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n887_), .A2(new_n429_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n654_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(G148gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n907_), .A2(new_n549_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  AND3_X1   g715(.A1(new_n907_), .A2(G162gat), .A3(new_n612_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G162gat), .B1(new_n907_), .B2(new_n610_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1347gat));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n884_), .A2(new_n264_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR4_X1   g721(.A1(new_n883_), .A2(new_n685_), .A3(new_n492_), .A4(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n923_), .B2(new_n290_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n873_), .A2(new_n610_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n925_), .A2(new_n861_), .B1(new_n880_), .B2(new_n879_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n549_), .B1(new_n926_), .B2(new_n874_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n684_), .B(new_n921_), .C1(new_n927_), .C2(new_n834_), .ZN(new_n928_));
  OAI211_X1 g727(.A(KEYINPUT62), .B(G169gat), .C1(new_n928_), .C2(new_n492_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n923_), .A2(new_n311_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n924_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n924_), .A2(new_n929_), .A3(KEYINPUT121), .A4(new_n930_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1348gat));
  NOR2_X1   g734(.A1(new_n928_), .A2(new_n654_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(G176gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n928_), .B2(new_n550_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n928_), .A2(new_n550_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n285_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n928_), .B2(new_n875_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n731_), .A2(new_n286_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n928_), .B2(new_n943_), .ZN(G1351gat));
  INV_X1    g743(.A(new_n429_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n883_), .A2(new_n264_), .A3(new_n945_), .A4(new_n685_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n946_), .A2(new_n947_), .A3(G197gat), .A4(new_n493_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n882_), .A2(new_n550_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n834_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n945_), .A2(new_n264_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n951_), .A2(new_n684_), .A3(new_n493_), .A4(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT124), .B1(new_n953_), .B2(new_n273_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT123), .B1(new_n953_), .B2(new_n273_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n948_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n948_), .B2(new_n954_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n951_), .A2(new_n684_), .A3(new_n952_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n654_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(new_n271_), .ZN(G1353gat));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n550_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963_));
  OR2_X1    g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  OR3_X1    g763(.A1(new_n962_), .A2(new_n963_), .A3(new_n964_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n963_), .B1(new_n962_), .B2(new_n964_), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT63), .B(G211gat), .Z(new_n967_));
  AOI22_X1  g766(.A1(new_n965_), .A2(new_n966_), .B1(new_n962_), .B2(new_n967_), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n946_), .B2(new_n610_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n612_), .A2(G218gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT126), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n969_), .B1(new_n946_), .B2(new_n971_), .ZN(G1355gat));
endmodule


