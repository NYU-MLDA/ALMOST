//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT22), .B(G169gat), .Z(new_n206_));
  OAI211_X1 g005(.A(new_n204_), .B(new_n205_), .C1(G176gat), .C2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n203_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT30), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  INV_X1    g019(.A(G113gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(G120gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n219_), .B(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G15gat), .B(G43gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT31), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G99gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n226_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT2), .ZN(new_n237_));
  OR2_X1    g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT3), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(KEYINPUT3), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT85), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT85), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT83), .Z(new_n245_));
  NAND2_X1  g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT84), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(KEYINPUT1), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(KEYINPUT1), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n238_), .A3(new_n236_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT29), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT88), .B(G197gat), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n257_), .B(KEYINPUT21), .C1(new_n258_), .C2(new_n256_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G211gat), .B(G218gat), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(G204gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n258_), .B2(G204gat), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n259_), .B(new_n261_), .C1(new_n263_), .C2(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT21), .A3(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(G228gat), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT87), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n254_), .A2(new_n266_), .B1(KEYINPUT89), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT89), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n254_), .A2(new_n266_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n272_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G22gat), .B(G50gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT28), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n253_), .A2(KEYINPUT29), .A3(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G78gat), .B(G106gat), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n279_), .B1(new_n253_), .B2(KEYINPUT29), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(KEYINPUT90), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n275_), .B(new_n286_), .C1(new_n272_), .C2(new_n271_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n280_), .A2(new_n283_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(KEYINPUT91), .ZN(new_n289_));
  OAI22_X1  g088(.A1(new_n276_), .A2(new_n284_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n287_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT92), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n289_), .A2(new_n287_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n284_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT92), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n297_), .B(new_n298_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n253_), .B(new_n223_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n253_), .A2(new_n305_), .A3(new_n223_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n303_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n306_), .B(new_n307_), .C1(new_n301_), .C2(new_n305_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G29gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT33), .ZN(new_n317_));
  XOR2_X1   g116(.A(G8gat), .B(G36gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(G64gat), .B(G92gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT19), .Z(new_n325_));
  XOR2_X1   g124(.A(new_n266_), .B(new_n217_), .Z(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(KEYINPUT20), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n266_), .B(new_n217_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n329_));
  INV_X1    g128(.A(new_n325_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n323_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(KEYINPUT20), .A3(new_n325_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n322_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n314_), .A2(new_n315_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n302_), .A2(new_n307_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n313_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n306_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n339_), .B(new_n340_), .C1(new_n341_), .C2(new_n307_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n317_), .A2(new_n336_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n304_), .A2(new_n308_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT96), .B1(new_n344_), .B2(new_n340_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n314_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n304_), .A2(new_n308_), .A3(KEYINPUT96), .A4(new_n313_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n334_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  OAI21_X1  g150(.A(new_n343_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n300_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n294_), .A2(new_n299_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT98), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n332_), .A2(new_n355_), .A3(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT97), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT97), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n332_), .A2(new_n358_), .A3(new_n335_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT27), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(KEYINPUT97), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n354_), .A2(new_n348_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n235_), .B1(new_n353_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n366_), .A3(new_n362_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT100), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n234_), .B1(new_n347_), .B2(new_n346_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n300_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n363_), .A2(KEYINPUT99), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n300_), .A2(new_n374_), .A3(new_n372_), .A4(new_n367_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT100), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n365_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G230gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT64), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT7), .ZN(new_n380_));
  INV_X1    g179(.A(G99gat), .ZN(new_n381_));
  INV_X1    g180(.A(G106gat), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .A4(KEYINPUT67), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384_));
  OAI22_X1  g183(.A1(new_n384_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G99gat), .A2(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n383_), .A2(new_n385_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G85gat), .B(G92gat), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT8), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT8), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G57gat), .A2(G64gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G57gat), .A2(G64gat), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(new_n399_), .A3(KEYINPUT11), .ZN(new_n400_));
  AND2_X1   g199(.A1(G71gat), .A2(G78gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G71gat), .A2(G78gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT68), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT11), .ZN(new_n405_));
  INV_X1    g204(.A(G57gat), .ZN(new_n406_));
  INV_X1    g205(.A(G64gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n408_), .B2(new_n397_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n405_), .A3(new_n397_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT68), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n401_), .A2(new_n402_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n404_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n411_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT10), .B(G99gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT65), .B1(new_n419_), .B2(G106gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT9), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT9), .B1(new_n425_), .B2(KEYINPUT66), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n388_), .A2(new_n389_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n381_), .A2(KEYINPUT10), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n381_), .A2(KEYINPUT10), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n382_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n420_), .A2(new_n427_), .A3(new_n429_), .A4(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n396_), .A2(new_n414_), .A3(new_n418_), .A4(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n418_), .A2(new_n414_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n390_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n394_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n440_), .A3(KEYINPUT12), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n379_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n379_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT69), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(KEYINPUT69), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G120gat), .B(G148gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n256_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT5), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(new_n212_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n455_), .A2(KEYINPUT70), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT70), .B1(new_n455_), .B2(new_n456_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n459_), .A2(KEYINPUT13), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(KEYINPUT13), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G1gat), .A2(G8gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT14), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G15gat), .A2(G22gat), .ZN(new_n465_));
  AND2_X1   g264(.A1(G15gat), .A2(G22gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G15gat), .B(G22gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(G1gat), .A2(G8gat), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(new_n463_), .A3(new_n471_), .A4(new_n464_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G50gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G43gat), .ZN(new_n475_));
  INV_X1    g274(.A(G43gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G50gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(G29gat), .A2(G36gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n477_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n473_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n483_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G29gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n484_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n469_), .A2(new_n472_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(new_n496_), .A3(KEYINPUT79), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n485_), .A2(new_n486_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT79), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n494_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT80), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n497_), .A2(KEYINPUT80), .A3(new_n502_), .A4(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n493_), .A2(KEYINPUT15), .A3(new_n495_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n494_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n498_), .A3(new_n487_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n511_), .A2(KEYINPUT81), .A3(new_n498_), .A4(new_n487_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n507_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT82), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n211_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n507_), .A2(new_n516_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n462_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n377_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n473_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(new_n436_), .Z(new_n530_));
  NOR2_X1   g329(.A1(new_n530_), .A2(KEYINPUT17), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G183gat), .B(G211gat), .Z(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  MUX2_X1   g335(.A(KEYINPUT17), .B(new_n531_), .S(new_n536_), .Z(new_n537_));
  NOR2_X1   g336(.A1(new_n530_), .A2(KEYINPUT77), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n537_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n439_), .A2(new_n500_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT34), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n509_), .A2(new_n510_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n439_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n439_), .B2(new_n500_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(new_n544_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n553_), .A3(new_n545_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n544_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n545_), .ZN(new_n557_));
  OAI221_X1 g356(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT36), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G134gat), .ZN(new_n562_));
  INV_X1    g361(.A(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n554_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n560_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n541_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n571_), .A2(KEYINPUT37), .A3(new_n567_), .A4(new_n565_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n540_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT78), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n527_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n575_), .A2(G1gat), .A3(new_n348_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT38), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT102), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(KEYINPUT38), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n526_), .B(KEYINPUT101), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n375_), .A2(KEYINPUT100), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n375_), .A2(KEYINPUT100), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n353_), .A2(new_n364_), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n581_), .A2(new_n582_), .B1(new_n583_), .B2(new_n235_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n568_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n571_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n540_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n580_), .A2(new_n584_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n348_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n579_), .A3(new_n590_), .ZN(G1324gat));
  INV_X1    g390(.A(new_n370_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(G8gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n575_), .A2(G8gat), .A3(new_n370_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(G8gat), .A3(new_n595_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n588_), .B2(new_n235_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT41), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n235_), .A2(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n575_), .B2(new_n606_), .ZN(G1326gat));
  OR3_X1    g406(.A1(new_n575_), .A2(G22gat), .A3(new_n300_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n588_), .A2(new_n354_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G22gat), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(KEYINPUT42), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT42), .B1(new_n611_), .B2(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(G1327gat));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n570_), .A2(new_n572_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n584_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n377_), .A2(KEYINPUT43), .A3(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n540_), .B(new_n580_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n348_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n584_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT43), .B1(new_n377_), .B2(new_n619_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n627_), .A2(KEYINPUT44), .A3(new_n540_), .A4(new_n580_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT105), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n623_), .A2(new_n631_), .A3(new_n624_), .A4(new_n628_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(G29gat), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n540_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n586_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n527_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n348_), .A2(G29gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT106), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT107), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n623_), .A2(new_n592_), .A3(new_n628_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G36gat), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n637_), .A2(KEYINPUT45), .A3(new_n646_), .A4(new_n592_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n527_), .A2(new_n646_), .A3(new_n636_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(new_n370_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n643_), .B1(new_n645_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n643_), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n651_), .C1(new_n644_), .C2(G36gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(G1329gat));
  NAND4_X1  g455(.A1(new_n623_), .A2(G43gat), .A3(new_n235_), .A4(new_n628_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n476_), .B1(new_n638_), .B2(new_n234_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g459(.A1(new_n623_), .A2(new_n354_), .A3(new_n628_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n623_), .A2(KEYINPUT108), .A3(new_n354_), .A4(new_n628_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(G50gat), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n637_), .A2(new_n474_), .A3(new_n354_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1331gat));
  NOR2_X1   g466(.A1(new_n377_), .A2(new_n525_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT110), .ZN(new_n669_));
  INV_X1    g468(.A(new_n462_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n574_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT109), .Z(new_n672_));
  AND2_X1   g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G57gat), .B1(new_n673_), .B2(new_n624_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n525_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n584_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n670_), .A2(new_n587_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(new_n406_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n624_), .B2(new_n678_), .ZN(G1332gat));
  NOR2_X1   g478(.A1(new_n676_), .A2(new_n677_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n407_), .B1(new_n680_), .B2(new_n592_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT48), .Z(new_n682_));
  NOR2_X1   g481(.A1(new_n370_), .A2(G64gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT111), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n673_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n680_), .B2(new_n235_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n673_), .A2(new_n687_), .A3(new_n235_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1334gat));
  INV_X1    g490(.A(G78gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n673_), .A2(new_n692_), .A3(new_n354_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n680_), .B2(new_n354_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(KEYINPUT50), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT50), .B1(new_n696_), .B2(new_n697_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n693_), .B1(new_n698_), .B2(new_n699_), .ZN(G1335gat));
  NOR3_X1   g499(.A1(new_n462_), .A2(new_n635_), .A3(new_n634_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n669_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n624_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n462_), .A2(new_n525_), .A3(new_n634_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n627_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(G85gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n624_), .B2(new_n707_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n703_), .B2(new_n592_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n706_), .A2(new_n592_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(G92gat), .B2(new_n710_), .ZN(G1337gat));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT114), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(new_n235_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G99gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n234_), .A2(new_n419_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n669_), .A2(new_n701_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n713_), .A2(KEYINPUT114), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n716_), .A2(new_n720_), .A3(new_n718_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(new_n714_), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n627_), .A2(new_n354_), .A3(new_n705_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n354_), .A2(new_n382_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n702_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  OAI221_X1 g529(.A(new_n730_), .B1(new_n702_), .B2(new_n727_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  NAND3_X1  g531(.A1(new_n441_), .A2(new_n379_), .A3(new_n443_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n441_), .A2(new_n443_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n445_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT55), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n444_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n734_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT56), .B1(new_n740_), .B2(new_n453_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n735_), .B2(new_n445_), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT55), .B(new_n379_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n733_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n454_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n741_), .A2(new_n525_), .A3(new_n456_), .A4(new_n746_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n497_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n511_), .A2(new_n499_), .A3(new_n487_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n521_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n524_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n524_), .A2(KEYINPUT116), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n748_), .B(new_n749_), .C1(new_n459_), .C2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT57), .A3(new_n635_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n757_), .A2(new_n456_), .A3(new_n746_), .A4(new_n741_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(KEYINPUT117), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n744_), .A2(new_n745_), .A3(new_n454_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n745_), .B1(new_n744_), .B2(new_n454_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n456_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n765_), .B1(new_n769_), .B2(new_n757_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n617_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n757_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n617_), .B(KEYINPUT118), .C1(new_n764_), .C2(new_n770_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n759_), .A2(new_n635_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n761_), .B1(new_n780_), .B2(KEYINPUT120), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n634_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n573_), .A2(new_n460_), .A3(new_n675_), .A4(new_n461_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n592_), .A2(new_n354_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n624_), .A3(new_n235_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT119), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n776_), .A2(new_n760_), .A3(new_n779_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n787_), .B1(new_n794_), .B2(new_n540_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n791_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(new_n221_), .A3(new_n675_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n798_), .ZN(new_n802_));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n525_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n800_), .B2(new_n462_), .ZN(new_n805_));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n462_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n802_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n806_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(G1341gat));
  INV_X1    g608(.A(G127gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n800_), .A2(new_n810_), .A3(new_n540_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G127gat), .B1(new_n802_), .B2(new_n634_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1342gat));
  INV_X1    g612(.A(G134gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n800_), .A2(new_n814_), .A3(new_n619_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G134gat), .B1(new_n802_), .B2(new_n586_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1343gat));
  NAND3_X1  g616(.A1(new_n370_), .A2(new_n354_), .A3(new_n234_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n795_), .A2(new_n348_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n525_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n670_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n634_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1346gat));
  AOI21_X1  g625(.A(G162gat), .B1(new_n819_), .B2(new_n586_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n617_), .A2(G162gat), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT121), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n819_), .B2(new_n829_), .ZN(G1347gat));
  NAND2_X1  g629(.A1(new_n592_), .A2(new_n372_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n354_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n525_), .B(new_n832_), .C1(new_n784_), .C2(new_n787_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n833_), .A2(new_n206_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT122), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n836_), .A2(new_n837_), .A3(new_n841_), .A4(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1348gat));
  AND2_X1   g642(.A1(new_n788_), .A2(new_n832_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G176gat), .B1(new_n844_), .B2(new_n670_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n795_), .A2(new_n354_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n831_), .A2(new_n462_), .A3(new_n212_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1349gat));
  NOR2_X1   g647(.A1(new_n831_), .A2(new_n540_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G183gat), .B1(new_n846_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n540_), .A2(new_n208_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n844_), .B2(new_n851_), .ZN(G1350gat));
  NAND2_X1  g651(.A1(new_n844_), .A2(new_n617_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G190gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n844_), .A2(new_n209_), .A3(new_n586_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1351gat));
  NAND2_X1  g655(.A1(new_n354_), .A2(new_n348_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n796_), .A2(new_n858_), .A3(new_n234_), .A4(new_n592_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n675_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT123), .B(G197gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1352gat));
  NOR2_X1   g661(.A1(new_n859_), .A2(new_n462_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n256_), .ZN(G1353gat));
  INV_X1    g663(.A(new_n859_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n540_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n869_), .A2(new_n870_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n870_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n868_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1354gat));
  OAI21_X1  g674(.A(KEYINPUT125), .B1(new_n859_), .B2(new_n635_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n795_), .A2(new_n857_), .A3(new_n235_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n592_), .A4(new_n586_), .ZN(new_n879_));
  INV_X1    g678(.A(G218gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n865_), .A2(G218gat), .A3(new_n617_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT126), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n882_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1355gat));
endmodule


