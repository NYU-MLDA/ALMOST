//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G22gat), .B(G50gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G78gat), .B(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G155gat), .ZN(new_n210_));
  INV_X1    g009(.A(G162gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT81), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G155gat), .B2(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n218_), .A2(new_n219_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n212_), .A2(new_n229_), .A3(new_n214_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n212_), .A2(new_n229_), .A3(new_n214_), .A4(KEYINPUT82), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(new_n233_), .C1(KEYINPUT1), .C2(new_n215_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G141gat), .B(G148gat), .Z(new_n235_));
  AND3_X1   g034(.A1(new_n234_), .A2(KEYINPUT83), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT83), .B1(new_n234_), .B2(new_n235_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n228_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT85), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(new_n228_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(KEYINPUT29), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n246_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(G197gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT87), .B1(new_n246_), .B2(G197gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT88), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT21), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT21), .B1(new_n248_), .B2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n252_), .B(new_n258_), .C1(new_n250_), .C2(KEYINPUT21), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G228gat), .ZN(new_n261_));
  INV_X1    g060(.A(G233gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n245_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n234_), .A2(new_n235_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n234_), .A2(KEYINPUT83), .A3(new_n235_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n271_), .B2(new_n228_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n260_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n263_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n244_), .B1(new_n265_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n244_), .A3(new_n274_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n209_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n279_), .A2(new_n275_), .A3(new_n208_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n203_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n208_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n277_), .A3(new_n209_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n202_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT92), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n292_), .B1(new_n294_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT94), .ZN(new_n302_));
  INV_X1    g101(.A(G183gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT23), .B1(new_n303_), .B2(new_n297_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT79), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n303_), .A2(new_n297_), .A3(KEYINPUT23), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n305_), .A2(new_n306_), .B1(new_n291_), .B2(new_n287_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT94), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n293_), .A2(KEYINPUT92), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n293_), .A2(KEYINPUT92), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n299_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n311_), .B2(new_n292_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT22), .B(G169gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n290_), .B1(new_n314_), .B2(new_n289_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n306_), .A2(new_n304_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n313_), .A2(new_n318_), .B1(new_n259_), .B2(new_n255_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n305_), .A2(new_n306_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n320_), .B2(new_n317_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n297_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n295_), .B2(G190gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n293_), .A2(new_n296_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT78), .ZN(new_n326_));
  NOR3_X1   g125(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n290_), .A2(new_n328_), .A3(new_n291_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n327_), .B(new_n329_), .C1(new_n306_), .C2(new_n304_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n321_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(new_n260_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n319_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT95), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n273_), .A2(new_n321_), .A3(new_n331_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n313_), .A2(new_n318_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT20), .B(new_n340_), .C1(new_n341_), .C2(new_n273_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n337_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n273_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n260_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT20), .A3(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(new_n337_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  INV_X1    g148(.A(G92gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT18), .B(G64gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n339_), .A2(new_n344_), .A3(new_n348_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(new_n337_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n353_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n358_), .A3(KEYINPUT27), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n339_), .A2(new_n348_), .A3(new_n344_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n355_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT101), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n359_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n242_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n271_), .A2(new_n228_), .A3(new_n377_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT4), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n374_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n380_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n374_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n373_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n373_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n382_), .A2(new_n386_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n391_), .A2(KEYINPUT4), .B1(new_n382_), .B2(new_n383_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n387_), .B(new_n390_), .C1(new_n392_), .C2(new_n374_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT99), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n387_), .B1(new_n392_), .B2(new_n374_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT99), .A3(new_n373_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n377_), .B(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT80), .B(G71gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT30), .B(G99gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G15gat), .B(G43gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT31), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n332_), .B(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n405_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR4_X1   g209(.A1(new_n286_), .A2(new_n368_), .A3(new_n399_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT98), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n379_), .A2(new_n412_), .A3(new_n380_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT98), .B1(new_n382_), .B2(new_n386_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(G225gat), .A4(G233gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n381_), .A2(new_n374_), .A3(new_n384_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n390_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n389_), .A2(KEYINPUT33), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n373_), .C1(new_n385_), .C2(new_n388_), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n417_), .B(new_n362_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n357_), .A2(KEYINPUT32), .A3(new_n354_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n339_), .A2(new_n344_), .A3(new_n348_), .A4(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n395_), .A2(new_n397_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n285_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT100), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT100), .B(new_n285_), .C1(new_n421_), .C2(new_n426_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n359_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n367_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n365_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n286_), .A2(new_n433_), .A3(new_n398_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n430_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n411_), .B1(new_n435_), .B2(new_n410_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G15gat), .B(G22gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(G1gat), .A2(G8gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(KEYINPUT14), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT73), .ZN(new_n440_));
  XOR2_X1   g239(.A(G1gat), .B(G8gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G43gat), .B(G50gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(G29gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT15), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT74), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n441_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n440_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450_));
  INV_X1    g249(.A(new_n446_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n445_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G229gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT75), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n447_), .A2(new_n452_), .A3(new_n454_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n449_), .A2(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G229gat), .A3(G233gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n458_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(G71gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT67), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G71gat), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n475_), .A2(new_n477_), .A3(G78gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(G78gat), .B1(new_n475_), .B2(new_n477_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G57gat), .A2(G64gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT11), .B1(new_n486_), .B2(new_n481_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT68), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(KEYINPUT11), .C1(new_n486_), .C2(new_n481_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n480_), .A2(new_n485_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n490_), .ZN(new_n492_));
  INV_X1    g291(.A(G78gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n476_), .A2(G71gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n474_), .A2(KEYINPUT67), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n475_), .A2(new_n477_), .A3(G78gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n485_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n491_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT10), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G99gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT64), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n504_), .A3(KEYINPUT64), .ZN(new_n507_));
  AOI21_X1  g306(.A(G106gat), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(G85gat), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n350_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n350_), .A2(G85gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(G92gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n510_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  INV_X1    g326(.A(G106gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n501_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(new_n522_), .A3(new_n523_), .A4(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n517_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n508_), .A2(new_n526_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n473_), .B1(new_n500_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n533_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n514_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n507_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n528_), .B1(new_n544_), .B2(new_n505_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n541_), .A2(new_n542_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n480_), .A2(new_n488_), .A3(new_n490_), .A4(new_n485_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n492_), .A2(new_n498_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n539_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n500_), .A2(KEYINPUT12), .A3(new_n536_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n541_), .A2(new_n542_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n543_), .A2(new_n545_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n552_), .B(new_n553_), .C1(new_n491_), .C2(new_n499_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n473_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n538_), .A2(new_n550_), .A3(new_n551_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n473_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n546_), .A2(new_n549_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT5), .B(G176gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n557_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n472_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n536_), .A2(new_n445_), .ZN(new_n580_));
  AOI211_X1 g379(.A(new_n579_), .B(new_n580_), .C1(new_n451_), .C2(new_n536_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n578_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT71), .Z(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n584_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n442_), .B(new_n500_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G211gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT16), .B(G183gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n601_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR4_X1   g409(.A1(new_n436_), .A2(new_n575_), .A3(new_n597_), .A4(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n398_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT103), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n436_), .A2(new_n575_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n596_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n585_), .A2(new_n590_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT37), .A3(new_n595_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n610_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n622_), .A2(G1gat), .A3(new_n398_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n623_), .A2(KEYINPUT104), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT104), .B1(new_n623_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n623_), .A2(new_n624_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n623_), .A2(new_n629_), .A3(new_n624_), .ZN(new_n630_));
  OAI221_X1 g429(.A(new_n614_), .B1(new_n625_), .B2(new_n626_), .C1(new_n628_), .C2(new_n630_), .ZN(G1324gat));
  NOR3_X1   g430(.A1(new_n622_), .A2(G8gat), .A3(new_n433_), .ZN(new_n632_));
  INV_X1    g431(.A(G8gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n611_), .B2(new_n368_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n632_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n638_), .B(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n611_), .B2(new_n409_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT41), .Z(new_n644_));
  NOR3_X1   g443(.A1(new_n622_), .A2(G15gat), .A3(new_n410_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  XNOR2_X1  g445(.A(new_n285_), .B(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G22gat), .B1(new_n612_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n648_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n622_), .B2(new_n651_), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n435_), .A2(new_n410_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n411_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n597_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n610_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n575_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n398_), .A2(G29gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT107), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n664_), .A3(new_n620_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n620_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n436_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n658_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n670_), .B(new_n659_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n669_), .A2(new_n671_), .A3(new_n398_), .ZN(new_n672_));
  INV_X1    g471(.A(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n663_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n669_), .A2(new_n671_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n368_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n660_), .A2(new_n676_), .A3(new_n368_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n675_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n679_), .B(KEYINPUT45), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n669_), .A2(new_n671_), .A3(new_n433_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n683_), .B(KEYINPUT46), .C1(new_n676_), .C2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1329gat));
  INV_X1    g485(.A(new_n669_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n658_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n687_), .A2(G43gat), .A3(new_n409_), .A4(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n656_), .A2(new_n410_), .A3(new_n659_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n690_), .A2(G43gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n660_), .B2(new_n647_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n286_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n677_), .B2(new_n698_), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n621_), .A2(new_n573_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n471_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n655_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n399_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n573_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n471_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n655_), .A2(new_n596_), .A3(new_n657_), .A4(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n398_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n706_), .A2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n709_), .B2(new_n433_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n433_), .A2(G64gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n704_), .B2(new_n715_), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n709_), .B2(new_n410_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT49), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n705_), .A2(new_n474_), .A3(new_n409_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  OAI21_X1  g519(.A(G78gat), .B1(new_n709_), .B2(new_n648_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT50), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n705_), .A2(new_n493_), .A3(new_n647_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n708_), .A2(new_n610_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n656_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n399_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n665_), .A2(new_n667_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n725_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n509_), .A2(G85gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n513_), .B1(new_n398_), .B2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n727_), .B1(new_n732_), .B2(new_n734_), .ZN(G1336gat));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n350_), .A3(new_n368_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n433_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n350_), .ZN(G1337gat));
  OAI211_X1 g537(.A(new_n726_), .B(new_n409_), .C1(new_n505_), .C2(new_n544_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n728_), .A2(new_n410_), .A3(new_n725_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n501_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n741_), .B(new_n742_), .Z(G1338gat));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n528_), .A3(new_n286_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n668_), .A2(new_n286_), .A3(new_n610_), .A4(new_n708_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  NAND4_X1  g552(.A1(new_n433_), .A2(new_n399_), .A3(new_n409_), .A4(new_n285_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT115), .Z(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n550_), .A2(new_n551_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n558_), .B1(new_n757_), .B2(new_n559_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n557_), .A2(new_n759_), .A3(KEYINPUT55), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT55), .B1(new_n557_), .B2(new_n759_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT69), .B(new_n558_), .C1(new_n546_), .C2(new_n549_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n555_), .B1(new_n554_), .B2(new_n473_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n757_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(KEYINPUT111), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n557_), .A2(new_n759_), .A3(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n758_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n763_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n756_), .B1(new_n773_), .B2(new_n566_), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT56), .B(new_n568_), .C1(new_n763_), .C2(new_n772_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n471_), .A4(new_n569_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n461_), .A2(new_n456_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n447_), .A2(new_n454_), .A3(new_n452_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n779_), .B(new_n467_), .C1(new_n456_), .C2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n470_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n570_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n771_), .B1(new_n770_), .B2(new_n758_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n758_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT112), .B(new_n786_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n566_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT56), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n756_), .B(new_n566_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n471_), .A3(new_n569_), .A4(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT113), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n778_), .A2(new_n784_), .A3(new_n792_), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT114), .B(KEYINPUT57), .C1(new_n793_), .C2(new_n596_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n596_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n776_), .A2(new_n569_), .A3(new_n782_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n569_), .A4(new_n782_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n620_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n794_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n793_), .A2(new_n596_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT114), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n657_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n621_), .A2(new_n472_), .A3(new_n707_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT54), .Z(new_n809_));
  OAI21_X1  g608(.A(new_n755_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT57), .B1(new_n793_), .B2(new_n596_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n610_), .B1(new_n801_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n808_), .B(KEYINPUT54), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n755_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT59), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n810_), .A2(KEYINPUT59), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n817_), .A2(G113gat), .A3(new_n471_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n795_), .A2(new_n800_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n803_), .A2(new_n821_), .A3(new_n804_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n806_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n809_), .B1(new_n823_), .B2(new_n610_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n819_), .B1(new_n824_), .B2(new_n815_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT116), .B(new_n755_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n471_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n818_), .A2(new_n828_), .ZN(G1340gat));
  XNOR2_X1  g628(.A(KEYINPUT117), .B(G120gat), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n817_), .B2(new_n573_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(KEYINPUT60), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n833_), .B(new_n835_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n832_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n816_), .A2(new_n814_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n822_), .A2(new_n795_), .A3(new_n800_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n811_), .A2(new_n821_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n610_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n815_), .B1(new_n841_), .B2(new_n813_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n830_), .B1(new_n844_), .B2(new_n707_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n827_), .A2(new_n834_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n845_), .B(new_n846_), .C1(new_n847_), .C2(new_n833_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n837_), .A2(new_n848_), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n827_), .B2(new_n657_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n657_), .A2(G127gat), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(KEYINPUT119), .Z(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n817_), .B2(new_n852_), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n841_), .A2(new_n813_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n855_), .B2(new_n755_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n819_), .B(new_n815_), .C1(new_n841_), .C2(new_n813_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n854_), .B(new_n597_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n620_), .B(new_n838_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G134gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n858_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n368_), .A2(new_n398_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n855_), .A2(new_n410_), .A3(new_n286_), .A4(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n472_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT121), .B(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n707_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n223_), .ZN(G1345gat));
  OAI21_X1  g670(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n610_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n824_), .A2(new_n409_), .A3(new_n285_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n657_), .A4(new_n865_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n872_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n866_), .A2(new_n211_), .A3(new_n666_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n873_), .A2(new_n597_), .A3(new_n865_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n211_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n433_), .A2(new_n399_), .A3(new_n410_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n814_), .A2(new_n648_), .A3(new_n885_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n288_), .B(new_n884_), .C1(new_n886_), .C2(new_n471_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n888_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n471_), .A3(new_n314_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n886_), .B2(new_n573_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n855_), .A2(KEYINPUT124), .A3(new_n285_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n824_), .B2(new_n286_), .ZN(new_n896_));
  AND4_X1   g695(.A1(new_n573_), .A2(new_n894_), .A3(new_n896_), .A4(new_n885_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n897_), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g697(.A(new_n886_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n899_), .A2(new_n294_), .A3(new_n610_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n894_), .A2(new_n896_), .A3(new_n657_), .A4(new_n885_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n303_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n899_), .B2(new_n666_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n886_), .A2(new_n300_), .A3(new_n597_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n433_), .A2(new_n399_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n873_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n472_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n256_), .ZN(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n707_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(new_n911_), .ZN(G1353gat));
  AND2_X1   g713(.A1(new_n873_), .A2(new_n906_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n657_), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n915_), .A2(new_n657_), .A3(new_n919_), .A4(new_n916_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1354gat));
  AOI21_X1  g722(.A(G218gat), .B1(new_n915_), .B2(new_n597_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n620_), .A2(G218gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT127), .Z(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n915_), .B2(new_n926_), .ZN(G1355gat));
endmodule


