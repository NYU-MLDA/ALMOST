//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  OR2_X1    g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n202_), .B(new_n203_), .C1(new_n206_), .C2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G113gat), .ZN(new_n214_));
  INV_X1    g013(.A(G120gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G113gat), .A2(G120gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n211_), .A2(new_n216_), .A3(new_n212_), .A4(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n225_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n202_), .A4(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n204_), .B(KEYINPUT88), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n207_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n210_), .A2(new_n221_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n210_), .A2(new_n229_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n219_), .A2(new_n232_), .A3(new_n220_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n232_), .B2(new_n220_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n230_), .A2(KEYINPUT99), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n231_), .A2(new_n234_), .A3(KEYINPUT99), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT100), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT4), .B1(new_n235_), .B2(new_n236_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n231_), .A2(new_n234_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT4), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n239_), .B1(new_n243_), .B2(new_n238_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G85gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(G1gat), .B(G29gat), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n244_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255_));
  INV_X1    g054(.A(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT83), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n263_));
  AND4_X1   g062(.A1(KEYINPUT83), .A2(new_n258_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G190gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT80), .B(G183gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G183gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT81), .B1(new_n271_), .B2(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n269_), .A3(G183gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n266_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n256_), .A2(new_n257_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT24), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n275_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n271_), .A2(KEYINPUT80), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n271_), .A2(KEYINPUT80), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT25), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n280_), .A2(new_n283_), .A3(KEYINPUT82), .A4(new_n267_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n265_), .A2(new_n276_), .A3(new_n279_), .A4(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(G176gat), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT84), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n254_), .B1(G190gat), .B2(new_n268_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(KEYINPUT84), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n278_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT87), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(new_n234_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G227gat), .A2(G233gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  MUX2_X1   g101(.A(new_n220_), .B(new_n221_), .S(new_n232_), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n296_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n300_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n302_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n251_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT92), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT96), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G211gat), .B(G218gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n320_), .ZN(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(G204gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G197gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT21), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n327_), .A3(new_n319_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n317_), .B1(new_n293_), .B2(new_n330_), .ZN(new_n331_));
  AOI211_X1 g130(.A(KEYINPUT96), .B(new_n329_), .C1(new_n285_), .C2(new_n292_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT94), .B1(new_n286_), .B2(new_n287_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n257_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n278_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n286_), .A2(KEYINPUT94), .A3(new_n287_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n336_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n343_));
  AOI21_X1  g142(.A(G176gat), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n278_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT95), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n254_), .B1(G183gat), .B2(G190gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n254_), .A2(new_n258_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n267_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n349_), .B(new_n279_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n329_), .A3(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT20), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n316_), .B1(new_n333_), .B2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G8gat), .B(G36gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n348_), .A2(new_n354_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n330_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n285_), .A2(new_n292_), .A3(new_n329_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(KEYINPUT20), .A3(new_n316_), .A4(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n357_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n293_), .A2(new_n330_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT96), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n293_), .A2(new_n317_), .A3(new_n330_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n356_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n315_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n362_), .B1(new_n374_), .B2(new_n367_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n312_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n363_), .B1(new_n357_), .B2(new_n368_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n315_), .B1(new_n333_), .B2(new_n356_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n365_), .A2(KEYINPUT20), .ZN(new_n379_));
  INV_X1    g178(.A(new_n366_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n379_), .A2(new_n316_), .A3(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n377_), .B(KEYINPUT27), .C1(new_n382_), .C2(new_n363_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n376_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n210_), .A2(new_n385_), .A3(new_n229_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT28), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n386_), .B(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n330_), .ZN(new_n391_));
  INV_X1    g190(.A(G228gat), .ZN(new_n392_));
  INV_X1    g191(.A(G233gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n390_), .B(new_n330_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G78gat), .B(G106gat), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT90), .B(new_n389_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n399_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n389_), .A2(KEYINPUT90), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(new_n395_), .A3(new_n396_), .A4(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n397_), .A2(new_n399_), .A3(new_n389_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n384_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n311_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n309_), .A2(new_n310_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT98), .B1(new_n369_), .B2(new_n375_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n374_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n377_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n238_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n249_), .B1(new_n243_), .B2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n235_), .A2(new_n236_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT33), .B1(new_n244_), .B2(new_n249_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NOR4_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n239_), .A4(new_n248_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n415_), .A2(new_n418_), .A3(new_n422_), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n357_), .B2(new_n368_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n250_), .B(new_n430_), .C1(new_n382_), .C2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n410_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT101), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n384_), .A2(new_n251_), .A3(new_n409_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(KEYINPUT101), .A3(new_n410_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n412_), .B1(new_n414_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT75), .B(G1gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT76), .B(G8gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT14), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G15gat), .B(G22gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G1gat), .ZN(new_n446_));
  INV_X1    g245(.A(G1gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n448_));
  AOI21_X1  g247(.A(G8gat), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(G8gat), .A3(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G71gat), .B(G78gat), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n456_), .A3(KEYINPUT11), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G231gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n452_), .B(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G127gat), .B(G155gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(G183gat), .B(G211gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(KEYINPUT17), .B2(new_n467_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n462_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT65), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(KEYINPUT65), .ZN(new_n478_));
  OR2_X1    g277(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n479_), .A2(G92gat), .A3(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n476_), .B(new_n478_), .C1(new_n481_), .C2(KEYINPUT9), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n485_), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n488_), .A3(KEYINPUT66), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT7), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n483_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n501_), .A2(new_n493_), .A3(new_n488_), .A4(KEYINPUT66), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(new_n495_), .A3(new_n500_), .A4(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G85gat), .B(G92gat), .Z(new_n504_));
  AOI21_X1  g303(.A(new_n491_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n491_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n495_), .A2(new_n502_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n486_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n490_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT68), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n490_), .B(new_n511_), .C1(new_n505_), .C2(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n459_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n459_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n490_), .A2(KEYINPUT69), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n490_), .A2(KEYINPUT69), .ZN(new_n520_));
  OAI22_X1  g319(.A1(new_n519_), .A2(new_n520_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(KEYINPUT12), .A3(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G230gat), .A2(G233gat), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n516_), .A2(new_n518_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n514_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n513_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(G120gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n528_), .A3(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT72), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(KEYINPUT72), .A3(new_n538_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n474_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(KEYINPUT13), .A3(new_n543_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT73), .B(G43gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G50gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G29gat), .B(G36gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT79), .B1(new_n452_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT79), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n549_), .B(new_n550_), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n553_), .B(new_n554_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n555_));
  OAI22_X1  g354(.A1(new_n552_), .A2(new_n555_), .B1(new_n551_), .B2(new_n452_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n551_), .B(KEYINPUT15), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n451_), .A3(new_n450_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n561_), .B(new_n557_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n256_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n323_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n547_), .A2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n439_), .A2(new_n473_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n521_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n517_), .A2(new_n551_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n578_), .A2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G134gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(G162gat), .Z(new_n590_));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n590_), .B(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n594_), .A3(new_n586_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n574_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(new_n595_), .A3(new_n574_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n573_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n602_), .A2(new_n251_), .A3(new_n440_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n593_), .A2(new_n595_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n573_), .A2(KEYINPUT103), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n438_), .A2(new_n414_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n412_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n572_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n607_), .A3(new_n472_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n251_), .B1(new_n608_), .B2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n605_), .B1(new_n447_), .B2(new_n616_), .ZN(G1324gat));
  NOR2_X1   g416(.A1(new_n613_), .A2(new_n384_), .ZN(new_n618_));
  INV_X1    g417(.A(G8gat), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n621_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n384_), .A2(new_n441_), .ZN(new_n625_));
  OAI22_X1  g424(.A1(new_n623_), .A2(new_n624_), .B1(new_n602_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n601_), .A2(new_n629_), .A3(new_n413_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n608_), .A2(new_n615_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n413_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(new_n632_), .B2(G15gat), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n634_), .B(new_n629_), .C1(new_n631_), .C2(new_n413_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT104), .B(new_n630_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n601_), .A2(new_n641_), .A3(new_n409_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n631_), .B2(new_n409_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT101), .B1(new_n432_), .B2(new_n410_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n434_), .B(new_n409_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n413_), .B1(new_n652_), .B2(new_n436_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n649_), .B(new_n599_), .C1(new_n653_), .C2(new_n412_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT105), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n600_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n611_), .A2(new_n657_), .A3(new_n649_), .A4(new_n599_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n572_), .A2(new_n472_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(KEYINPUT44), .A3(new_n660_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n250_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G29gat), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n611_), .A2(new_n606_), .A3(new_n660_), .ZN(new_n667_));
  INV_X1    g466(.A(G29gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n250_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n648_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT106), .B(new_n671_), .C1(new_n665_), .C2(G29gat), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1328gat));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n384_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n667_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n659_), .A2(KEYINPUT44), .A3(new_n660_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT44), .B1(new_n659_), .B2(new_n660_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n384_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n680_), .B2(new_n674_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT46), .B(new_n677_), .C1(new_n680_), .C2(new_n674_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1329gat));
  AND4_X1   g484(.A1(G43gat), .A2(new_n663_), .A3(new_n413_), .A4(new_n664_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G43gat), .B1(new_n667_), .B2(new_n413_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT47), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n678_), .A2(new_n679_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(G43gat), .A3(new_n413_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  INV_X1    g490(.A(new_n687_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n667_), .B2(new_n409_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n409_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n689_), .B2(new_n696_), .ZN(G1331gat));
  INV_X1    g496(.A(new_n547_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n593_), .A2(new_n595_), .A3(new_n574_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n570_), .A2(new_n472_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n596_), .A3(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n611_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n250_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT107), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n547_), .A2(new_n571_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n606_), .A2(new_n473_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n611_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(G57gat), .A3(new_n250_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n704_), .A2(new_n709_), .ZN(G1332gat));
  INV_X1    g509(.A(new_n702_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n711_), .A2(G64gat), .A3(new_n384_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G64gat), .B1(new_n707_), .B2(new_n384_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(KEYINPUT48), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT48), .B1(new_n714_), .B2(new_n715_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n712_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT109), .B(new_n712_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n707_), .B2(new_n414_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT110), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n711_), .A2(G71gat), .A3(new_n414_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  OR3_X1    g526(.A1(new_n711_), .A2(G78gat), .A3(new_n410_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G78gat), .B1(new_n707_), .B2(new_n410_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT111), .Z(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT50), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT50), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n705_), .A2(new_n473_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n439_), .A2(new_n734_), .A3(new_n607_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n250_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n734_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n659_), .A2(new_n737_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n250_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n735_), .B2(new_n675_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n675_), .A2(G92gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n742_), .ZN(G1337gat));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n659_), .A2(new_n413_), .A3(new_n737_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G99gat), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n413_), .A2(new_n487_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n735_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n747_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n746_), .B2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n744_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n753_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(KEYINPUT51), .A3(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n735_), .A2(new_n488_), .A3(new_n409_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n659_), .A2(new_n409_), .A3(new_n737_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G106gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n758_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  OAI21_X1  g566(.A(new_n538_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n524_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n524_), .B2(new_n770_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n516_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n525_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n769_), .B1(new_n776_), .B2(new_n535_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n773_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n775_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n524_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n536_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n768_), .B1(new_n777_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n556_), .A2(new_n557_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n561_), .B(new_n558_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n565_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n567_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT57), .B(new_n607_), .C1(new_n783_), .C2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n538_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n569_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n567_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n776_), .A2(new_n769_), .A3(new_n535_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n536_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n788_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n607_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n791_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n607_), .B1(new_n783_), .B2(new_n788_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n787_), .A2(new_n792_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT58), .B(new_n805_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n599_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n804_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n473_), .B1(new_n801_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n547_), .A2(new_n701_), .A3(new_n814_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n413_), .A2(new_n384_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n818_), .A2(new_n250_), .A3(new_n410_), .A4(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n214_), .B1(new_n821_), .B2(new_n570_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT117), .Z(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT118), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n825_), .B(KEYINPUT59), .C1(KEYINPUT118), .C2(new_n821_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n570_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n828_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g628(.A(new_n821_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n215_), .B1(new_n547_), .B2(KEYINPUT60), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT120), .Z(new_n832_));
  OAI211_X1 g631(.A(new_n830_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n215_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n547_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n215_), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n830_), .B2(new_n472_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n473_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n830_), .B2(new_n606_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n600_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n413_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n842_), .A2(new_n250_), .A3(new_n409_), .A4(new_n384_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n570_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT122), .B(G141gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n846_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT123), .B(G148gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n850_), .A2(new_n698_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n850_), .B2(new_n698_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1345gat));
  AOI21_X1  g653(.A(new_n473_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n855_), .B(new_n857_), .ZN(G1346gat));
  AOI21_X1  g657(.A(G162gat), .B1(new_n850_), .B2(new_n606_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n600_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(G162gat), .B2(new_n860_), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n311_), .A2(new_n384_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n818_), .A2(new_n571_), .A3(new_n410_), .A4(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n409_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(KEYINPUT125), .A3(new_n571_), .A4(new_n862_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(G169gat), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n866_), .A2(new_n862_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n571_), .C1(new_n338_), .C2(new_n337_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n865_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n867_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n870_), .A2(KEYINPUT126), .A3(new_n872_), .A4(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1348gat));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(G176gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n871_), .A2(new_n698_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(G176gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n881_), .B2(new_n880_), .ZN(G1349gat));
  INV_X1    g683(.A(new_n871_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n473_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n268_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n886_), .B2(new_n352_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n885_), .B2(new_n600_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n871_), .A2(new_n606_), .A3(new_n267_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  AND2_X1   g690(.A1(new_n842_), .A2(new_n409_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n384_), .A2(new_n250_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n570_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n323_), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n547_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n325_), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n892_), .A2(new_n472_), .A3(new_n893_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n899_), .B2(new_n900_), .ZN(G1354gat));
  NOR2_X1   g702(.A1(new_n894_), .A2(new_n607_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(G218gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n894_), .A2(new_n600_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(G218gat), .B2(new_n906_), .ZN(G1355gat));
endmodule


