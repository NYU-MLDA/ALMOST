//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203_));
  INV_X1    g002(.A(G120gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G113gat), .ZN(new_n205_));
  INV_X1    g004(.A(G113gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(new_n214_), .B2(KEYINPUT25), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n213_), .A2(new_n215_), .A3(new_n217_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n221_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT83), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G183gat), .A3(G190gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT23), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(G183gat), .B2(G190gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G169gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI22_X1  g045(.A1(new_n231_), .A2(new_n239_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G99gat), .ZN(new_n248_));
  INV_X1    g047(.A(G43gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(G15gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT30), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT31), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n251_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n212_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n209_), .A2(new_n211_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n267_));
  INV_X1    g066(.A(G155gat), .ZN(new_n268_));
  INV_X1    g067(.A(G162gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT85), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(G155gat), .B2(G162gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275_));
  INV_X1    g074(.A(G141gat), .ZN(new_n276_));
  INV_X1    g075(.A(G148gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n273_), .A2(KEYINPUT1), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G155gat), .A3(G162gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n270_), .A2(new_n286_), .A3(new_n272_), .A4(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G141gat), .B(G148gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n263_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n212_), .A2(new_n285_), .A3(new_n291_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT93), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n297_), .A3(KEYINPUT4), .A4(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(new_n293_), .B2(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT95), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n293_), .A2(new_n294_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n300_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n305_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT33), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n302_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n300_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n310_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT95), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n314_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n304_), .A2(KEYINPUT33), .A3(new_n313_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n293_), .A2(KEYINPUT4), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(new_n301_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n299_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n310_), .B1(new_n312_), .B2(new_n301_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT19), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT89), .ZN(new_n329_));
  AND2_X1   g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n329_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT21), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT88), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT89), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n332_), .A2(KEYINPUT21), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n334_), .A2(new_n341_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT20), .B1(new_n247_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n240_), .A2(new_n242_), .ZN(new_n349_));
  INV_X1    g148(.A(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT26), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n218_), .A2(G183gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n215_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n223_), .A2(new_n221_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n349_), .A2(new_n227_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n236_), .A2(new_n238_), .B1(G183gat), .B2(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n245_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n357_), .A2(new_n359_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n328_), .B1(new_n348_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n247_), .A2(new_n347_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n357_), .A2(new_n359_), .A3(new_n344_), .A4(new_n346_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n328_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n362_), .A2(KEYINPUT20), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n372_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G64gat), .B(G92gat), .Z(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n378_), .B2(new_n370_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n368_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n372_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n367_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n366_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n361_), .A2(new_n384_), .A3(new_n365_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n321_), .A2(new_n326_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n267_), .B1(new_n320_), .B2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n314_), .A2(new_n319_), .A3(new_n315_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n316_), .A2(new_n318_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n391_), .A2(KEYINPUT33), .B1(new_n324_), .B2(new_n325_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n361_), .A2(new_n384_), .A3(new_n365_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n384_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n390_), .A2(new_n392_), .A3(KEYINPUT96), .A4(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n361_), .A2(new_n365_), .A3(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n348_), .A2(new_n328_), .A3(new_n360_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n227_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n401_), .A2(new_n349_), .B1(new_n358_), .B2(new_n245_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT89), .B1(new_n339_), .B2(new_n340_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n343_), .B1(new_n340_), .B2(new_n335_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n345_), .B1(new_n405_), .B2(new_n341_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n400_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n364_), .B1(new_n407_), .B2(new_n362_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n399_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n310_), .B1(new_n304_), .B2(new_n317_), .ZN(new_n410_));
  OAI221_X1 g209(.A(new_n398_), .B1(new_n409_), .B2(new_n397_), .C1(new_n410_), .C2(new_n391_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n389_), .A2(new_n396_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G22gat), .B(G50gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT28), .B1(new_n292_), .B2(KEYINPUT29), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n292_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n413_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT90), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n292_), .B2(KEYINPUT29), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n347_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT86), .ZN(new_n430_));
  INV_X1    g229(.A(G228gat), .ZN(new_n431_));
  INV_X1    g230(.A(G233gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n434_), .A3(new_n347_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n433_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n425_), .B(new_n426_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n417_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n424_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n440_), .B(new_n436_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n412_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n439_), .A2(new_n444_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n410_), .A2(new_n391_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n380_), .A2(KEYINPUT97), .A3(new_n383_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT97), .B1(new_n380_), .B2(new_n383_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(new_n399_), .B2(new_n408_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n387_), .A3(KEYINPUT27), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .A4(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n266_), .B1(new_n446_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n261_), .A2(new_n264_), .A3(new_n448_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n450_), .A2(new_n459_), .A3(new_n455_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n445_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT99), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT99), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n464_), .B(new_n445_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n457_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G85gat), .B(G92gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT10), .B(G99gat), .Z(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT6), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT9), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n470_), .A2(new_n473_), .A3(new_n475_), .A4(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(G99gat), .B(G106gat), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n484_), .A3(new_n475_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n468_), .B(KEYINPUT66), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT8), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(KEYINPUT8), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n479_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G29gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT34), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n494_), .B(new_n479_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n496_), .A2(KEYINPUT74), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n500_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n496_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n501_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n496_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT76), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G134gat), .B(G162gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT36), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(KEYINPUT36), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n512_), .A2(new_n518_), .B1(new_n519_), .B2(new_n510_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n467_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G230gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT68), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(KEYINPUT11), .B2(new_n524_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n491_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n491_), .A2(new_n531_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n523_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT69), .ZN(new_n535_));
  INV_X1    g334(.A(new_n532_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(KEYINPUT70), .A3(new_n530_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(KEYINPUT12), .A4(new_n491_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n491_), .A2(new_n538_), .A3(KEYINPUT12), .A4(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT71), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n536_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT12), .B1(new_n491_), .B2(new_n531_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n523_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n535_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT5), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G176gat), .B(G204gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT73), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n535_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT77), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n494_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n495_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n494_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G169gat), .B(G197gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT80), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n578_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n570_), .B(new_n585_), .Z(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(new_n531_), .Z(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT79), .ZN(new_n589_));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n540_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n594_), .B1(new_n597_), .B2(new_n586_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n586_), .B2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n561_), .A2(new_n584_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n522_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n448_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n202_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n467_), .A2(new_n583_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n516_), .B(KEYINPUT75), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n510_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n510_), .A2(new_n519_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n520_), .A2(KEYINPUT37), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n561_), .A2(new_n612_), .A3(new_n600_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n607_), .A2(new_n613_), .A3(new_n202_), .A4(new_n604_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n605_), .B1(new_n606_), .B2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n606_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT101), .ZN(G1324gat));
  NOR2_X1   g420(.A1(new_n460_), .A2(new_n461_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n565_), .B1(new_n603_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT39), .Z(new_n624_));
  NAND4_X1  g423(.A1(new_n607_), .A2(new_n613_), .A3(new_n565_), .A4(new_n622_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1325gat));
  NAND2_X1  g427(.A1(new_n607_), .A2(new_n613_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(G15gat), .A3(new_n265_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT102), .Z(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n602_), .B2(new_n265_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n633_), .A3(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n602_), .B2(new_n445_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n445_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n629_), .B2(new_n639_), .ZN(G1327gat));
  OAI211_X1 g439(.A(new_n583_), .B(new_n600_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n612_), .B1(new_n457_), .B2(new_n466_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  OAI221_X1 g444(.A(new_n612_), .B1(KEYINPUT104), .B2(new_n645_), .C1(new_n457_), .C2(new_n466_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT105), .B1(new_n647_), .B2(KEYINPUT44), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n646_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n641_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(G29gat), .A3(new_n604_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n560_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n600_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n521_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n607_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n448_), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n650_), .A2(new_n656_), .B1(G29gat), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT106), .ZN(G1328gat));
  OR2_X1    g464(.A1(new_n622_), .A2(KEYINPUT107), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n622_), .A2(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n662_), .A2(G36gat), .A3(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT45), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n651_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n647_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n622_), .A3(new_n655_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1329gat));
  XOR2_X1   g480(.A(KEYINPUT110), .B(G43gat), .Z(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n662_), .B2(new_n265_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n265_), .A2(new_n249_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n647_), .B2(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n684_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n687_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT112), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n650_), .B2(new_n685_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n691_), .A4(new_n683_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n693_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1330gat));
  NAND3_X1  g499(.A1(new_n676_), .A2(new_n447_), .A3(new_n655_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT113), .B1(new_n701_), .B2(G50gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n445_), .A2(G50gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT114), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n702_), .A2(new_n703_), .B1(new_n662_), .B2(new_n705_), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n659_), .A2(new_n583_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n467_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n612_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n660_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n604_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n659_), .A2(new_n583_), .A3(new_n600_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n522_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(G57gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n604_), .B2(KEYINPUT115), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(KEYINPUT115), .B2(new_n715_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n711_), .B1(new_n714_), .B2(new_n717_), .ZN(G1332gat));
  OAI21_X1  g517(.A(G64gat), .B1(new_n713_), .B2(new_n669_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT117), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n710_), .A2(new_n723_), .A3(new_n668_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n713_), .B2(new_n265_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT49), .ZN(new_n727_));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n710_), .A2(new_n728_), .A3(new_n266_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n713_), .B2(new_n445_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n710_), .A2(new_n733_), .A3(new_n447_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  NAND2_X1  g534(.A1(new_n708_), .A2(new_n661_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n476_), .B1(new_n736_), .B2(new_n448_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n651_), .A2(new_n600_), .A3(new_n707_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n448_), .A2(new_n476_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT118), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT119), .Z(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n739_), .B2(new_n669_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n736_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n477_), .A3(new_n622_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1337gat));
  NAND2_X1  g546(.A1(new_n266_), .A2(new_n471_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n736_), .A2(new_n748_), .B1(KEYINPUT120), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n738_), .A2(new_n266_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(G99gat), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(KEYINPUT120), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n752_), .B(new_n753_), .Z(G1338gat));
  AOI21_X1  g553(.A(new_n472_), .B1(new_n738_), .B2(new_n447_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT52), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n472_), .A3(new_n447_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n558_), .A2(new_n583_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT121), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n558_), .A2(KEYINPUT121), .A3(new_n583_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n523_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n549_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n545_), .A2(KEYINPUT55), .A3(new_n523_), .A4(new_n548_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n555_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n555_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n767_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n556_), .A2(new_n558_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n581_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n578_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n571_), .A2(new_n572_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n575_), .A2(new_n576_), .A3(new_n573_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT122), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT122), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n778_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n521_), .B1(new_n777_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n558_), .A2(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT123), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n558_), .A2(KEYINPUT123), .A3(new_n786_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n555_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n555_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n774_), .B(new_n796_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n709_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n794_), .B(KEYINPUT58), .C1(new_n795_), .C2(new_n797_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n788_), .A2(new_n789_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT57), .B(new_n521_), .C1(new_n777_), .C2(new_n787_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n660_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n613_), .A2(new_n584_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n448_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n265_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n206_), .A3(new_n583_), .A4(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n805_), .B(KEYINPUT54), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n802_), .A2(new_n803_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n660_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT59), .A3(new_n604_), .A4(new_n810_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n604_), .B(new_n810_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n584_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n811_), .B1(new_n819_), .B2(new_n206_), .ZN(G1340gat));
  OAI21_X1  g619(.A(new_n204_), .B1(new_n659_), .B2(KEYINPUT60), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n204_), .A2(KEYINPUT60), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n809_), .A2(new_n810_), .A3(new_n821_), .A4(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n659_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n204_), .ZN(G1341gat));
  INV_X1    g624(.A(G127gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n816_), .B2(new_n600_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT124), .B(new_n826_), .C1(new_n816_), .C2(new_n600_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n815_), .A2(new_n818_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n600_), .A2(new_n826_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n829_), .A2(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n809_), .A2(new_n834_), .A3(new_n520_), .A4(new_n810_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n709_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1343gat));
  NOR3_X1   g636(.A1(new_n668_), .A2(new_n445_), .A3(new_n266_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n809_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G141gat), .B1(new_n839_), .B2(new_n584_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n809_), .A2(new_n276_), .A3(new_n583_), .A4(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1344gat));
  OAI21_X1  g641(.A(G148gat), .B1(new_n839_), .B2(new_n659_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n809_), .A2(new_n277_), .A3(new_n561_), .A4(new_n838_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1345gat));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n839_), .B2(new_n600_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n809_), .A2(new_n660_), .A3(new_n838_), .A4(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n839_), .B2(new_n709_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n809_), .A2(new_n269_), .A3(new_n520_), .A4(new_n838_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  NOR3_X1   g652(.A1(new_n669_), .A2(new_n447_), .A3(new_n458_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n583_), .B(new_n854_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT62), .B1(new_n855_), .B2(KEYINPUT22), .ZN(new_n856_));
  OAI21_X1  g655(.A(G169gat), .B1(new_n855_), .B2(KEYINPUT62), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G169gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n856_), .ZN(G1348gat));
  INV_X1    g659(.A(new_n854_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n808_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n561_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g663(.A1(new_n808_), .A2(new_n600_), .A3(new_n861_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(G183gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n354_), .A2(new_n215_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n868_), .B2(new_n865_), .ZN(G1350gat));
  NAND3_X1  g668(.A1(new_n862_), .A2(new_n213_), .A3(new_n520_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n814_), .A2(new_n612_), .A3(new_n854_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(G190gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n871_), .B2(G190gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n870_), .B1(new_n873_), .B2(new_n874_), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n447_), .A2(new_n448_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n669_), .A2(new_n876_), .A3(new_n266_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n814_), .A2(new_n583_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(G197gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT126), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n808_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n882_), .A2(new_n883_), .A3(G197gat), .A4(new_n583_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n879_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n880_), .A2(new_n884_), .A3(new_n885_), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n561_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g687(.A(KEYINPUT63), .B(G211gat), .Z(new_n889_));
  NAND4_X1  g688(.A1(new_n814_), .A2(new_n660_), .A3(new_n877_), .A4(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n660_), .B(new_n877_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n892_), .A2(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n882_), .A2(new_n898_), .A3(new_n520_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n808_), .A2(new_n709_), .A3(new_n881_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(G1355gat));
endmodule


