//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT68), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT69), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT7), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n217_));
  OAI211_X1 g016(.A(G99gat), .B(G106gat), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n215_), .A2(new_n218_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(new_n203_), .B(new_n205_), .C1(new_n224_), .C2(new_n229_), .ZN(new_n230_));
  AND4_X1   g029(.A1(KEYINPUT70), .A2(new_n224_), .A3(KEYINPUT8), .A4(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n202_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n227_), .B2(KEYINPUT9), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT66), .B(G92gat), .Z(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(new_n225_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n233_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT64), .B(G106gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT10), .B(G99gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n222_), .A2(new_n218_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n224_), .A2(new_n229_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n203_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n204_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n224_), .A2(KEYINPUT70), .A3(KEYINPUT8), .A4(new_n229_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT72), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n232_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G71gat), .B(G78gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(KEYINPUT11), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT71), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253_));
  XOR2_X1   g052(.A(G57gat), .B(G64gat), .Z(new_n254_));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n252_), .A2(new_n257_), .B1(new_n255_), .B2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(KEYINPUT71), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n253_), .A3(new_n249_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT11), .A4(new_n250_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n262_), .A2(KEYINPUT12), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n248_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n245_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT12), .B1(new_n265_), .B2(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n269_), .B1(new_n273_), .B2(new_n267_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT5), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G176gat), .B(G204gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n279_), .B(KEYINPUT73), .Z(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n282_), .A2(KEYINPUT74), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n282_), .B2(new_n284_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G29gat), .B(G36gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT76), .ZN(new_n295_));
  INV_X1    g094(.A(G36gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G29gat), .ZN(new_n297_));
  INV_X1    g096(.A(G29gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G36gat), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT76), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT77), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n294_), .A2(KEYINPUT76), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G43gat), .B(G50gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n309_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n301_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G1gat), .ZN(new_n314_));
  INV_X1    g113(.A(G8gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT14), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G22gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G15gat), .ZN(new_n318_));
  INV_X1    g117(.A(G15gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G22gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(KEYINPUT81), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(KEYINPUT81), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G8gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n327_), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n313_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n310_), .A2(new_n326_), .A3(new_n312_), .A4(new_n328_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n312_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n311_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT15), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT15), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n310_), .A2(new_n339_), .A3(new_n312_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n329_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n330_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n335_), .B1(new_n344_), .B2(new_n331_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G141gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G169gat), .B(G197gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT85), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n345_), .A2(KEYINPUT86), .A3(new_n348_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n313_), .A2(new_n329_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n334_), .B1(new_n354_), .B2(new_n332_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n348_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n352_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n350_), .B1(new_n351_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n293_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT94), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(KEYINPUT94), .B2(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n366_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n370_), .A2(KEYINPUT94), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n368_), .A2(KEYINPUT2), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT3), .Z(new_n374_));
  OAI211_X1 g173(.A(new_n362_), .B(new_n364_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n362_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(KEYINPUT1), .B2(new_n362_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n373_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n365_), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G127gat), .B(G134gat), .Z(new_n381_));
  XOR2_X1   g180(.A(G113gat), .B(G120gat), .Z(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT91), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n382_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(KEYINPUT91), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n385_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT99), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT100), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n380_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n380_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT100), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n388_), .A2(KEYINPUT4), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n361_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT0), .ZN(new_n402_));
  INV_X1    g201(.A(G57gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(new_n225_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n361_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n400_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n405_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n399_), .B2(new_n407_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  INV_X1    g211(.A(G197gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(G204gat), .ZN(new_n414_));
  INV_X1    g213(.A(G204gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(G197gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT21), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n414_), .A2(KEYINPUT96), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT97), .B1(new_n415_), .B2(G197gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(KEYINPUT96), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n417_), .B(new_n418_), .C1(new_n424_), .C2(KEYINPUT21), .ZN(new_n425_));
  INV_X1    g224(.A(new_n418_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(KEYINPUT21), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(G169gat), .B2(G176gat), .ZN(new_n430_));
  NOR3_X1   g229(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT23), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT26), .B(G190gat), .Z(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT25), .B(G183gat), .Z(new_n436_));
  OAI211_X1 g235(.A(new_n432_), .B(new_n434_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(G183gat), .B2(G190gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT88), .B(G176gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G169gat), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n439_), .A2(new_n440_), .B1(G169gat), .B2(G176gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n428_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n425_), .A2(new_n427_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT87), .B(G183gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(KEYINPUT25), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n432_), .B(new_n434_), .C1(new_n448_), .C2(new_n435_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n434_), .B1(G190gat), .B2(new_n447_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(KEYINPUT89), .B2(new_n441_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n441_), .A2(KEYINPUT89), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n444_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n443_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n445_), .A2(new_n453_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G226gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT19), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  MUX2_X1   g261(.A(new_n456_), .B(new_n459_), .S(new_n462_), .Z(new_n463_));
  XNOR2_X1  g262(.A(G8gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT18), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n461_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n444_), .A2(KEYINPUT20), .A3(new_n462_), .A4(new_n454_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT103), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n463_), .A2(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n412_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n470_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n467_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(new_n412_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n409_), .B(new_n411_), .C1(new_n475_), .C2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT105), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n380_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n483_), .B(KEYINPUT28), .Z(new_n484_));
  XOR2_X1   g283(.A(G22gat), .B(G50gat), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n428_), .A2(KEYINPUT95), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n380_), .B2(new_n482_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G228gat), .A3(G233gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n487_), .B(new_n490_), .C1(new_n380_), .C2(new_n482_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT98), .Z(new_n493_));
  AND3_X1   g292(.A1(new_n489_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n491_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n489_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n485_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n484_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n501_), .A3(new_n484_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n453_), .B(KEYINPUT30), .ZN(new_n507_));
  XOR2_X1   g306(.A(G71gat), .B(G99gat), .Z(new_n508_));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G15gat), .B(G43gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT90), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n510_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n387_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n517_), .A2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n506_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n506_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n480_), .A2(new_n481_), .A3(new_n505_), .A4(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n496_), .A2(new_n501_), .A3(new_n484_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n528_), .B2(new_n502_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT105), .B1(new_n529_), .B2(new_n479_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n502_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n532_), .B2(new_n479_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n411_), .A2(new_n534_), .ZN(new_n535_));
  OAI221_X1 g334(.A(new_n410_), .B1(KEYINPUT101), .B2(KEYINPUT33), .C1(new_n399_), .C2(new_n407_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n406_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n361_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n405_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n477_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n409_), .A2(new_n411_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n476_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n463_), .B2(new_n542_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n505_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n533_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n533_), .B2(new_n546_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n531_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G190gat), .B(G218gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n271_), .A2(new_n313_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n248_), .A2(new_n561_), .A3(new_n341_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n248_), .B2(new_n341_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n559_), .A2(new_n556_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI221_X1 g365(.A(new_n560_), .B1(new_n556_), .B2(new_n559_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n555_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n553_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT79), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT80), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n566_), .A2(new_n567_), .A3(new_n574_), .A4(new_n571_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n568_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  AOI211_X1 g377(.A(new_n578_), .B(new_n568_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT83), .ZN(new_n584_));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT84), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT82), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n262_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n342_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n342_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n589_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n594_), .A3(new_n588_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n586_), .A2(new_n587_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n581_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n360_), .A2(new_n550_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n541_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n604_), .A2(G1gat), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT107), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n527_), .A2(new_n530_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n533_), .A2(new_n546_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT104), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n533_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n610_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n609_), .B1(new_n614_), .B2(new_n576_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n576_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n550_), .A2(KEYINPUT107), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n602_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n290_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n359_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n605_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n608_), .A2(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(new_n604_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n475_), .A2(new_n478_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n315_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n615_), .A2(new_n617_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(new_n620_), .A3(new_n625_), .A4(new_n601_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n629_), .B2(G8gat), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n627_), .A3(G8gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n626_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT40), .B(new_n626_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(new_n526_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n621_), .B2(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT41), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT41), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n624_), .A2(new_n319_), .A3(new_n526_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(G1326gat));
  NAND3_X1  g444(.A1(new_n624_), .A2(new_n317_), .A3(new_n532_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G22gat), .B1(new_n621_), .B2(new_n505_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(new_n620_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n576_), .A2(new_n602_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n614_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n541_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n614_), .A2(KEYINPUT43), .A3(new_n580_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n550_), .B2(new_n581_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n620_), .B(new_n602_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n614_), .B2(new_n580_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n550_), .A2(new_n656_), .A3(new_n581_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n601_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n660_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n605_), .A2(new_n298_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n654_), .B1(new_n665_), .B2(new_n666_), .ZN(G1328gat));
  NAND3_X1  g466(.A1(new_n653_), .A2(new_n296_), .A3(new_n625_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n669_));
  XOR2_X1   g468(.A(new_n668_), .B(new_n669_), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n660_), .A2(new_n664_), .A3(new_n625_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(G36gat), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT46), .ZN(G1329gat));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n640_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n660_), .A2(new_n664_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT110), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n660_), .A2(new_n664_), .A3(new_n678_), .A4(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n653_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(new_n640_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n685_), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  NAND4_X1  g486(.A1(new_n660_), .A2(new_n664_), .A3(G50gat), .A4(new_n532_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n681_), .A2(new_n505_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(G50gat), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT111), .Z(G1331gat));
  INV_X1    g490(.A(new_n293_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n358_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n618_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n541_), .A2(new_n696_), .A3(G57gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n696_), .B2(G57gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n581_), .A2(new_n290_), .A3(new_n602_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT112), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n614_), .A2(new_n358_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(KEYINPUT112), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n403_), .B1(new_n704_), .B2(new_n605_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n699_), .A2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT114), .Z(G1332gat));
  INV_X1    g506(.A(new_n625_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n704_), .A2(G64gat), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G64gat), .B1(new_n694_), .B2(new_n708_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT48), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT48), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1333gat));
  OR3_X1    g512(.A1(new_n704_), .A2(G71gat), .A3(new_n640_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n695_), .A2(new_n526_), .ZN(new_n715_));
  XOR2_X1   g514(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n715_), .A2(G71gat), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n715_), .B2(G71gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(G1334gat));
  OR3_X1    g519(.A1(new_n704_), .A2(G78gat), .A3(new_n505_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G78gat), .B1(new_n694_), .B2(new_n505_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT50), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT50), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1335gat));
  NOR2_X1   g524(.A1(new_n290_), .A2(new_n358_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n663_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n663_), .A2(KEYINPUT116), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n729_), .A2(KEYINPUT117), .A3(new_n730_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n541_), .A3(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n692_), .A2(new_n652_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n702_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n541_), .A2(new_n225_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n735_), .A2(new_n225_), .B1(new_n737_), .B2(new_n738_), .ZN(G1336gat));
  NOR2_X1   g538(.A1(new_n708_), .A2(new_n234_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n734_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n226_), .B1(new_n737_), .B2(new_n708_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OR3_X1    g542(.A1(new_n737_), .A2(new_n239_), .A3(new_n640_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n640_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n206_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g546(.A1(new_n737_), .A2(new_n238_), .A3(new_n505_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G106gat), .B1(new_n727_), .B2(new_n505_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT52), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT52), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n748_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NOR4_X1   g555(.A1(new_n288_), .A2(new_n289_), .A3(new_n358_), .A4(new_n602_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n580_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(new_n580_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n354_), .A2(new_n332_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n330_), .A2(new_n333_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n356_), .B1(new_n763_), .B2(new_n331_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n281_), .B(new_n765_), .C1(new_n351_), .C2(new_n357_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n264_), .A2(new_n268_), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n248_), .A2(new_n263_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n269_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n270_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n283_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n283_), .C1(new_n773_), .C2(new_n776_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n767_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n767_), .B(KEYINPUT58), .C1(new_n779_), .C2(new_n781_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n784_), .B(new_n785_), .C1(new_n577_), .C2(new_n579_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT86), .B1(new_n345_), .B2(new_n348_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n355_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n282_), .B1(new_n790_), .B2(new_n350_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n788_), .A2(new_n789_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n285_), .A2(new_n287_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n795_), .B2(new_n616_), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT57), .B(new_n576_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n786_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n761_), .B1(new_n602_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n605_), .A2(new_n625_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n799_), .A2(KEYINPUT59), .A3(new_n529_), .A4(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n358_), .A2(new_n281_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n777_), .A2(new_n778_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n780_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n778_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n794_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n616_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n795_), .A2(new_n787_), .A3(new_n616_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT119), .B1(new_n813_), .B2(new_n786_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n786_), .B(KEYINPUT119), .C1(new_n796_), .C2(new_n797_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n602_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n761_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n803_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n798_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n601_), .B1(new_n821_), .B2(new_n815_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(KEYINPUT120), .A3(new_n761_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n801_), .A2(new_n529_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n359_), .B(new_n802_), .C1(new_n826_), .C2(KEYINPUT59), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n358_), .A2(new_n828_), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n827_), .A2(new_n828_), .B1(new_n826_), .B2(new_n829_), .ZN(G1340gat));
  AOI211_X1 g629(.A(new_n692_), .B(new_n802_), .C1(new_n826_), .C2(KEYINPUT59), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n290_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n831_), .A2(new_n832_), .B1(new_n826_), .B2(new_n834_), .ZN(G1341gat));
  AOI211_X1 g634(.A(new_n602_), .B(new_n802_), .C1(new_n826_), .C2(KEYINPUT59), .ZN(new_n836_));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n601_), .A2(new_n837_), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n836_), .A2(new_n837_), .B1(new_n826_), .B2(new_n838_), .ZN(G1342gat));
  NAND2_X1  g638(.A1(new_n581_), .A2(G134gat), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n802_), .B(new_n840_), .C1(new_n826_), .C2(KEYINPUT59), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n824_), .A2(new_n576_), .A3(new_n825_), .ZN(new_n842_));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n842_), .A2(KEYINPUT121), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT121), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n841_), .A2(new_n844_), .A3(new_n845_), .ZN(G1343gat));
  NAND3_X1  g645(.A1(new_n817_), .A2(new_n818_), .A3(new_n803_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n822_), .B2(new_n761_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n505_), .A2(new_n526_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(new_n800_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n358_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n293_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n851_), .B2(new_n601_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n850_), .A2(new_n800_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n859_), .A2(KEYINPUT122), .A3(new_n602_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n856_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n851_), .A2(new_n857_), .A3(new_n601_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n859_), .B2(new_n602_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n856_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n851_), .B2(new_n576_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n581_), .A2(G162gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT123), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n851_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n708_), .A2(new_n541_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n526_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n505_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n799_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n359_), .ZN(new_n877_));
  INV_X1    g676(.A(G169gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(KEYINPUT62), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n440_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  OAI21_X1  g682(.A(new_n439_), .B1(new_n876_), .B2(new_n290_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT124), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n819_), .A2(new_n823_), .A3(new_n532_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n293_), .A2(G176gat), .A3(new_n873_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  AND3_X1   g687(.A1(new_n875_), .A2(new_n436_), .A3(new_n601_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n601_), .A3(new_n873_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n447_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n876_), .B2(new_n580_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n616_), .A2(new_n435_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT125), .Z(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n876_), .B2(new_n895_), .ZN(G1351gat));
  NAND4_X1  g695(.A1(new_n824_), .A2(KEYINPUT126), .A3(new_n849_), .A4(new_n871_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .A4(new_n871_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n359_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n413_), .ZN(G1352gat));
  AOI21_X1  g701(.A(new_n692_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n415_), .ZN(G1353gat));
  AOI21_X1  g703(.A(new_n602_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  NAND2_X1  g708(.A1(new_n581_), .A2(G218gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n616_), .B1(new_n897_), .B2(new_n900_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913_));
  AOI21_X1  g712(.A(G218gat), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n898_), .A2(new_n899_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n898_), .A2(new_n899_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n576_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT127), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n911_), .B1(new_n914_), .B2(new_n918_), .ZN(G1355gat));
endmodule


