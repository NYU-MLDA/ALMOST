//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  INV_X1    g000(.A(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT82), .B1(new_n203_), .B2(KEYINPUT22), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G169gat), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n202_), .B(new_n204_), .C1(new_n205_), .C2(KEYINPUT82), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n206_), .A2(new_n207_), .A3(new_n216_), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n214_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(KEYINPUT25), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT26), .B1(new_n214_), .B2(KEYINPUT80), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n223_));
  OAI21_X1  g022(.A(G183gat), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(G183gat), .C1(new_n222_), .C2(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n221_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n209_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT81), .B1(new_n208_), .B2(KEYINPUT23), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n211_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  MUX2_X1   g033(.A(new_n233_), .B(KEYINPUT24), .S(new_n234_), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n217_), .B1(new_n228_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G134gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G127gat), .ZN(new_n244_));
  INV_X1    g043(.A(G127gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G134gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT83), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT83), .B1(new_n244_), .B2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n246_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n247_), .A3(new_n241_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n240_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(G15gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n256_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT27), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n266_), .A2(G197gat), .ZN(new_n267_));
  INV_X1    g066(.A(G197gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(G204gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT21), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT90), .B1(new_n266_), .B2(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT90), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n268_), .A3(G204gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n274_), .C1(new_n268_), .C2(G204gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n270_), .B(new_n271_), .C1(new_n275_), .C2(KEYINPUT21), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT21), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n276_), .A2(new_n278_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n232_), .A2(new_n215_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n205_), .A2(new_n202_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n207_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT25), .B(G183gat), .Z(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT26), .B(G190gat), .Z(new_n286_));
  OAI211_X1 g085(.A(new_n235_), .B(new_n212_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n265_), .B1(new_n280_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n237_), .A2(new_n279_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n265_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT20), .A4(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n289_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n263_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT99), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT99), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n302_), .B(new_n263_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  INV_X1    g104(.A(G228gat), .ZN(new_n306_));
  INV_X1    g105(.A(G233gat), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT88), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(KEYINPUT88), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT89), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G155gat), .B(G162gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(KEYINPUT2), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT84), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT85), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n319_), .A2(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(KEYINPUT2), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G141gat), .ZN(new_n327_));
  INV_X1    g126(.A(G148gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT3), .ZN(new_n330_));
  OR3_X1    g129(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT86), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .A4(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n315_), .B1(new_n326_), .B2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n314_), .A2(KEYINPUT1), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n339_), .A3(new_n316_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n313_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n312_), .B1(new_n343_), .B2(new_n281_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n343_), .A2(new_n312_), .A3(new_n281_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n305_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n305_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G22gat), .B(G50gat), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n318_), .A2(new_n320_), .A3(KEYINPUT85), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n323_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n336_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n314_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n341_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n354_), .B1(new_n360_), .B2(new_n313_), .ZN(new_n361_));
  NOR4_X1   g160(.A1(new_n359_), .A2(KEYINPUT29), .A3(new_n341_), .A4(new_n353_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OR3_X1    g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n348_), .A2(KEYINPUT91), .A3(new_n344_), .A4(new_n349_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n352_), .A2(new_n365_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n366_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n347_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT92), .B(new_n305_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .A4(new_n350_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n255_), .B1(new_n359_), .B2(new_n341_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n337_), .A2(new_n254_), .A3(new_n250_), .A4(new_n342_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(KEYINPUT4), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT93), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n337_), .A2(new_n342_), .B1(new_n254_), .B2(new_n250_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G85gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT0), .B(G57gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT95), .B1(new_n384_), .B2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n385_), .A2(new_n389_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n377_), .A2(new_n383_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n385_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n389_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(KEYINPUT96), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n375_), .A2(new_n376_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n401_), .A2(new_n378_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n402_), .B2(new_n389_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n399_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n298_), .A2(new_n263_), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n280_), .A2(new_n288_), .A3(new_n265_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n265_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n297_), .B(KEYINPUT98), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n406_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n304_), .A2(new_n374_), .A3(new_n405_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n289_), .A2(new_n293_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n404_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n381_), .A2(new_n382_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n377_), .A2(new_n419_), .A3(new_n378_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n375_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n398_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n420_), .A2(KEYINPUT94), .A3(new_n398_), .A4(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n298_), .A2(new_n299_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n384_), .B2(new_n390_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n392_), .A2(KEYINPUT33), .A3(new_n394_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n374_), .B1(new_n418_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n413_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT97), .B(new_n374_), .C1(new_n418_), .C2(new_n431_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n262_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n304_), .A2(new_n412_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n374_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n262_), .A2(new_n404_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G22gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n258_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G15gat), .A2(G22gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G1gat), .A2(G8gat), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n447_), .A2(new_n448_), .B1(KEYINPUT14), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n445_), .B(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G43gat), .B(G50gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(G29gat), .B(G36gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G29gat), .B(G36gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n451_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT77), .Z(new_n464_));
  INV_X1    g263(.A(KEYINPUT15), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n458_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n455_), .A2(new_n456_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n452_), .A2(new_n453_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT15), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n451_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n473_), .A2(KEYINPUT76), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT76), .B1(new_n473_), .B2(new_n474_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n462_), .B(new_n464_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n451_), .B(new_n461_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G229gat), .A3(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT13), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT67), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G78gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT11), .ZN(new_n491_));
  INV_X1    g290(.A(new_n490_), .ZN(new_n492_));
  INV_X1    g291(.A(G64gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G57gat), .ZN(new_n494_));
  INV_X1    g293(.A(G57gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G64gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n496_), .A3(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n491_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510_));
  INV_X1    g309(.A(G99gat), .ZN(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n504_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n507_), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n514_), .B(new_n513_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n504_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G92gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT9), .ZN(new_n525_));
  AND2_X1   g324(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n501_), .A2(KEYINPUT9), .A3(new_n502_), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n512_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n506_), .A2(new_n508_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n500_), .B1(new_n523_), .B2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT65), .ZN(new_n536_));
  INV_X1    g335(.A(new_n514_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI211_X1 g338(.A(KEYINPUT8), .B(new_n503_), .C1(new_n539_), .C2(new_n533_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n521_), .B1(new_n520_), .B2(new_n504_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n500_), .B(new_n534_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(KEYINPUT65), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n542_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(KEYINPUT12), .B2(new_n535_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n534_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n500_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI211_X1 g354(.A(KEYINPUT66), .B(KEYINPUT12), .C1(new_n551_), .C2(new_n552_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n549_), .B(new_n545_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n547_), .B2(new_n557_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n488_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT36), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n459_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT15), .B1(new_n470_), .B2(new_n471_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n551_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT71), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n534_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n461_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n581_), .A2(new_n586_), .B1(new_n580_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n580_), .A2(new_n591_), .A3(new_n589_), .A4(new_n586_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n585_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n577_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n580_), .A2(new_n589_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n473_), .B2(new_n551_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n586_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n593_), .A4(new_n592_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n576_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n602_));
  INV_X1    g401(.A(new_n594_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n599_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n601_), .A2(KEYINPUT73), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n600_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n575_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT37), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n602_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n603_), .A2(new_n575_), .A3(new_n599_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(KEYINPUT37), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n620_), .B(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n500_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n474_), .B(new_n626_), .ZN(new_n627_));
  MUX2_X1   g426(.A(new_n623_), .B(new_n624_), .S(new_n627_), .Z(new_n628_));
  NAND2_X1  g427(.A1(new_n615_), .A2(new_n628_), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n442_), .A2(new_n486_), .A3(new_n571_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(G1gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n404_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n606_), .A2(KEYINPUT73), .A3(new_n575_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n611_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n601_), .A2(KEYINPUT73), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n442_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n486_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n570_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n628_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n405_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n634_), .A2(new_n635_), .A3(new_n646_), .ZN(G1324gat));
  XNOR2_X1  g446(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n648_));
  OAI21_X1  g447(.A(G8gat), .B1(new_n645_), .B2(new_n438_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(G8gat), .C1(new_n645_), .C2(new_n438_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(G8gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n630_), .A2(new_n654_), .A3(new_n437_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n648_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n648_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n655_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n657_), .B(new_n658_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n659_), .ZN(G1325gat));
  INV_X1    g459(.A(new_n645_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n262_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n258_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n630_), .A2(new_n258_), .A3(new_n662_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT102), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(G1326gat));
  OAI21_X1  g468(.A(G22gat), .B1(new_n645_), .B2(new_n439_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n630_), .A2(new_n446_), .A3(new_n374_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT37), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n613_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n436_), .A2(new_n441_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n610_), .A2(KEYINPUT103), .A3(new_n614_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n676_), .B2(new_n613_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n680_), .B1(new_n686_), .B2(KEYINPUT43), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n642_), .A2(new_n628_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n674_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n678_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n688_), .C1(new_n691_), .C2(new_n680_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G29gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n405_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n639_), .A2(new_n643_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n571_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n681_), .A2(new_n641_), .A3(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(new_n405_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n693_), .A2(new_n695_), .B1(new_n694_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT46), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n690_), .A2(new_n437_), .A3(new_n692_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n438_), .A2(G36gat), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n681_), .A2(new_n641_), .A3(new_n697_), .A4(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT45), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT45), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n707_), .A2(new_n708_), .B1(new_n701_), .B2(KEYINPUT46), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n704_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n702_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n712_), .B(new_n709_), .C1(new_n703_), .C2(G36gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1329gat));
  NAND4_X1  g513(.A1(new_n690_), .A2(G43gat), .A3(new_n662_), .A4(new_n692_), .ZN(new_n715_));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n698_), .B2(new_n262_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n720_), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  OR3_X1    g521(.A1(new_n698_), .A2(G50gat), .A3(new_n439_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n690_), .A2(new_n374_), .A3(new_n692_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n724_), .B2(G50gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NOR4_X1   g526(.A1(new_n442_), .A2(new_n641_), .A3(new_n570_), .A4(new_n629_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n495_), .A3(new_n404_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n639_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n485_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(new_n628_), .A3(new_n483_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n570_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n681_), .A2(new_n730_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n681_), .A2(KEYINPUT106), .A3(new_n730_), .A4(new_n733_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n404_), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n729_), .B1(new_n738_), .B2(new_n495_), .ZN(G1332gat));
  NAND2_X1  g538(.A1(new_n437_), .A2(new_n493_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT107), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n728_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n437_), .A3(new_n737_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G64gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n728_), .A2(new_n748_), .A3(new_n662_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n736_), .A2(new_n662_), .A3(new_n737_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT108), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n728_), .A2(new_n759_), .A3(new_n374_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n736_), .A2(new_n374_), .A3(new_n737_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(G78gat), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G78gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT110), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n696_), .A2(new_n570_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n681_), .A2(new_n486_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT111), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n681_), .A2(new_n773_), .A3(new_n486_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n404_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n570_), .A2(new_n641_), .A3(new_n628_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n779_));
  INV_X1    g578(.A(new_n680_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(KEYINPUT112), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n691_), .B2(new_n680_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n526_), .A2(new_n527_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n405_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n776_), .B1(new_n784_), .B2(new_n786_), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n524_), .B1(new_n784_), .B2(new_n437_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n775_), .A2(new_n524_), .A3(new_n437_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n438_), .B(new_n778_), .C1(new_n781_), .C2(new_n783_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT113), .B(new_n790_), .C1(new_n793_), .C2(new_n524_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1337gat));
  NAND2_X1  g594(.A1(new_n784_), .A2(new_n662_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G99gat), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n530_), .A2(new_n531_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n262_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n775_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  INV_X1    g601(.A(new_n800_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n802_), .B(new_n803_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n797_), .A2(new_n798_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n511_), .B1(new_n784_), .B2(new_n662_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n801_), .A2(new_n804_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(G1338gat));
  NAND3_X1  g609(.A1(new_n775_), .A2(new_n512_), .A3(new_n374_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n374_), .B(new_n777_), .C1(new_n691_), .C2(new_n680_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT52), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n512_), .B1(new_n813_), .B2(KEYINPUT52), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n812_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n811_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n486_), .A2(new_n825_), .A3(new_n628_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n732_), .A2(KEYINPUT116), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n570_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n615_), .A2(new_n824_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n615_), .B2(new_n828_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n464_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n462_), .B(new_n833_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n482_), .B1(new_n478_), .B2(new_n464_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n483_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n567_), .B2(new_n563_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n554_), .B1(new_n588_), .B2(new_n500_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT66), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n553_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n545_), .B1(new_n845_), .B2(new_n549_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n557_), .A2(KEYINPUT117), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(KEYINPUT55), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n557_), .A2(KEYINPUT117), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n562_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n841_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n845_), .A2(new_n549_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n546_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n542_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n859_), .B2(new_n545_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n855_), .B1(new_n860_), .B2(new_n849_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n557_), .A2(KEYINPUT117), .A3(new_n849_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT56), .B(new_n561_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n839_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n849_), .B1(new_n557_), .B2(KEYINPUT117), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n865_), .A3(new_n846_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n840_), .C1(new_n866_), .C2(new_n562_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n853_), .A2(new_n864_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n486_), .A2(new_n564_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n838_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n832_), .B1(new_n870_), .B2(new_n639_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n869_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n847_), .A2(KEYINPUT55), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n850_), .A3(new_n855_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n852_), .B1(new_n874_), .B2(new_n561_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n875_), .A2(new_n840_), .B1(new_n863_), .B2(new_n839_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n872_), .B1(new_n876_), .B2(new_n853_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n730_), .C1(new_n877_), .C2(new_n838_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n837_), .A2(new_n564_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n851_), .A2(KEYINPUT56), .ZN(new_n880_));
  INV_X1    g679(.A(new_n863_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(KEYINPUT58), .B(new_n879_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n677_), .A3(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n878_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n831_), .B1(new_n887_), .B2(new_n643_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n437_), .A2(new_n262_), .A3(new_n374_), .A4(new_n405_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n888_), .A2(new_n486_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n823_), .B1(new_n891_), .B2(G113gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n887_), .A2(new_n643_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n831_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n641_), .A3(new_n889_), .ZN(new_n896_));
  INV_X1    g695(.A(G113gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(KEYINPUT120), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n892_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT59), .B1(new_n895_), .B2(new_n889_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n888_), .A2(new_n902_), .A3(new_n890_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n895_), .A2(KEYINPUT59), .A3(new_n889_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(KEYINPUT121), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n486_), .A2(new_n897_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n899_), .B1(new_n908_), .B2(new_n909_), .ZN(G1340gat));
  NOR2_X1   g709(.A1(new_n888_), .A2(new_n890_), .ZN(new_n911_));
  INV_X1    g710(.A(G120gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n570_), .B2(KEYINPUT60), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(new_n913_), .C1(KEYINPUT60), .C2(new_n912_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n570_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n912_), .ZN(G1341gat));
  AOI21_X1  g715(.A(G127gat), .B1(new_n911_), .B2(new_n628_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n643_), .A2(new_n245_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n908_), .B2(new_n918_), .ZN(G1342gat));
  AOI21_X1  g718(.A(G134gat), .B1(new_n911_), .B2(new_n639_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n615_), .A2(new_n243_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n908_), .B2(new_n921_), .ZN(G1343gat));
  NOR3_X1   g721(.A1(new_n439_), .A2(new_n662_), .A3(new_n405_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n895_), .A2(new_n438_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n486_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n327_), .ZN(G1344gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n570_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n328_), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n924_), .A2(new_n643_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  INV_X1    g730(.A(G162gat), .ZN(new_n932_));
  NOR4_X1   g731(.A1(new_n924_), .A2(new_n932_), .A3(new_n684_), .A4(new_n682_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n924_), .B2(new_n730_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT122), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n936_), .B(new_n932_), .C1(new_n924_), .C2(new_n730_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n935_), .B2(new_n937_), .ZN(G1347gat));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n437_), .A2(new_n440_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n895_), .A2(new_n439_), .A3(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n486_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n939_), .B1(new_n943_), .B2(new_n203_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n205_), .ZN(new_n945_));
  OAI211_X1 g744(.A(KEYINPUT62), .B(G169gat), .C1(new_n942_), .C2(new_n486_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(G1348gat));
  OR3_X1    g746(.A1(new_n888_), .A2(KEYINPUT123), .A3(new_n374_), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT123), .B1(new_n888_), .B2(new_n374_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n940_), .A2(new_n202_), .A3(new_n570_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n202_), .B1(new_n942_), .B2(new_n570_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1349gat));
  NAND4_X1  g752(.A1(new_n948_), .A2(new_n628_), .A3(new_n941_), .A4(new_n949_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n942_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n628_), .A2(new_n285_), .ZN(new_n956_));
  AOI22_X1  g755(.A1(new_n954_), .A2(new_n213_), .B1(new_n955_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n942_), .B2(new_n615_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n730_), .A2(new_n286_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n942_), .B2(new_n959_), .ZN(G1351gat));
  NAND3_X1  g759(.A1(new_n405_), .A2(new_n374_), .A3(new_n262_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n888_), .A2(new_n438_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n486_), .B1(KEYINPUT124), .B2(new_n268_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n268_), .A2(KEYINPUT124), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(KEYINPUT125), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n964_), .B(new_n966_), .ZN(G1352gat));
  AND2_X1   g766(.A1(new_n962_), .A2(new_n571_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n266_), .A2(KEYINPUT126), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n266_), .A2(KEYINPUT126), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n968_), .B1(new_n969_), .B2(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n971_), .B1(new_n968_), .B2(new_n970_), .ZN(G1353gat));
  AOI211_X1 g771(.A(KEYINPUT63), .B(G211gat), .C1(new_n962_), .C2(new_n628_), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n962_), .A2(new_n628_), .ZN(new_n974_));
  XOR2_X1   g773(.A(KEYINPUT63), .B(G211gat), .Z(new_n975_));
  AOI21_X1  g774(.A(new_n973_), .B1(new_n974_), .B2(new_n975_), .ZN(G1354gat));
  INV_X1    g775(.A(G218gat), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n962_), .A2(new_n977_), .A3(new_n639_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n962_), .A2(new_n677_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n979_), .B2(new_n977_), .ZN(G1355gat));
endmodule


