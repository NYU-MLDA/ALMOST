//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT10), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT10), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G99gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AOI22_X1  g010(.A1(new_n206_), .A2(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n213_), .A2(G85gat), .A3(G92gat), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n218_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n215_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n206_), .A2(new_n207_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n209_), .A2(new_n211_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n215_), .A4(new_n220_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n202_), .A3(new_n207_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n227_), .A2(new_n230_), .A3(new_n202_), .A4(new_n207_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n218_), .A2(new_n219_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n221_), .B(new_n226_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G50gat), .ZN(new_n239_));
  INV_X1    g038(.A(G29gat), .ZN(new_n240_));
  INV_X1    g039(.A(G36gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G29gat), .A2(G36gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n239_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G50gat), .A3(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n238_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n226_), .A2(new_n221_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT68), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n232_), .A2(new_n234_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n255_), .B1(new_n256_), .B2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT15), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT15), .B1(new_n248_), .B2(new_n250_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT71), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT68), .B1(new_n235_), .B2(new_n236_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n254_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n265_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n253_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G232gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT34), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(KEYINPUT35), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n262_), .A2(KEYINPUT71), .A3(new_n266_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n271_), .B1(new_n270_), .B2(new_n265_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(KEYINPUT35), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n275_), .A2(KEYINPUT35), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .A4(new_n253_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G134gat), .ZN(new_n286_));
  INV_X1    g085(.A(G162gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n276_), .A2(new_n277_), .A3(new_n283_), .A4(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n276_), .A2(new_n283_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT36), .A3(new_n289_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n294_), .A2(KEYINPUT37), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT37), .B1(new_n294_), .B2(new_n296_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT13), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G57gat), .B(G64gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n304_));
  XOR2_X1   g103(.A(G71gat), .B(G78gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n303_), .A2(KEYINPUT11), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n237_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n238_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT67), .B1(new_n238_), .B2(new_n310_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n302_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G176gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G204gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n262_), .A2(KEYINPUT12), .A3(new_n308_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AND4_X1   g122(.A1(KEYINPUT70), .A2(new_n309_), .A3(new_n321_), .A4(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n237_), .B2(new_n308_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT70), .B1(new_n325_), .B2(new_n321_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n320_), .B(new_n311_), .C1(new_n324_), .C2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n315_), .B(new_n319_), .C1(new_n327_), .C2(new_n302_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n309_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(KEYINPUT70), .A3(new_n321_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(new_n301_), .A3(new_n320_), .A4(new_n311_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n319_), .B1(new_n335_), .B2(new_n315_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n300_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n315_), .B1(new_n327_), .B2(new_n302_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n319_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT13), .A3(new_n328_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G8gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT14), .ZN(new_n344_));
  AND2_X1   g143(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n347_), .B2(G1gat), .ZN(new_n348_));
  INV_X1    g147(.A(G15gat), .ZN(new_n349_));
  INV_X1    g148(.A(G22gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G15gat), .A2(G22gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n348_), .A2(G1gat), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G1gat), .ZN(new_n356_));
  OR2_X1    g155(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(G1gat), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT14), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n356_), .B1(new_n360_), .B2(new_n353_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n343_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(G1gat), .B1(new_n348_), .B2(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(G8gat), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(new_n252_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n251_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(G229gat), .A2(G233gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n368_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n366_), .B2(new_n265_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G141gat), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G197gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n373_), .B(new_n383_), .C1(new_n371_), .C2(new_n375_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n342_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT78), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n401_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n395_), .A2(new_n400_), .A3(new_n404_), .A4(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n378_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n378_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n393_), .A2(new_n394_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n408_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n409_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT81), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n408_), .A2(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT30), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n416_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G15gat), .B(G43gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n426_), .B(new_n429_), .Z(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n423_), .A3(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n426_), .B(new_n429_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n432_), .B(KEYINPUT81), .C1(new_n418_), .C2(new_n417_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(KEYINPUT83), .A3(new_n433_), .ZN(new_n437_));
  INV_X1    g236(.A(G120gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G127gat), .B(G134gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n439_), .A2(G113gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(G113gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n439_), .A2(G113gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(G113gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(G120gat), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n436_), .A2(new_n437_), .A3(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n437_), .A2(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G211gat), .B(G218gat), .Z(new_n452_));
  INV_X1    g251(.A(G204gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n380_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(KEYINPUT87), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G204gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n458_), .B2(new_n380_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n452_), .B1(new_n459_), .B2(KEYINPUT21), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT87), .B(G204gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT88), .B1(new_n461_), .B2(new_n380_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n463_), .A3(G197gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT21), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n380_), .A2(G204gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT21), .A3(new_n452_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G155gat), .B(G162gat), .Z(new_n472_));
  NAND2_X1  g271(.A1(G141gat), .A2(G148gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT85), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT2), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(KEYINPUT85), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT84), .A3(new_n482_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n476_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n472_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G155gat), .ZN(new_n487_));
  OR3_X1    g286(.A1(new_n487_), .A2(new_n287_), .A3(KEYINPUT1), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n287_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT1), .B1(new_n487_), .B2(new_n287_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n481_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(new_n473_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n486_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G78gat), .B(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  AND3_X1   g298(.A1(new_n471_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n471_), .B2(new_n496_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G22gat), .B(G50gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n486_), .A2(new_n504_), .A3(new_n494_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT28), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n474_), .A2(KEYINPUT2), .B1(new_n476_), .B2(KEYINPUT3), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n508_), .A2(new_n479_), .A3(new_n484_), .A4(new_n483_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n509_), .A2(new_n472_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(new_n504_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(KEYINPUT28), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n507_), .A3(new_n504_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n503_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n502_), .A2(KEYINPUT86), .A3(new_n512_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n471_), .A2(new_n496_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n499_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n471_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT86), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n516_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n517_), .A2(KEYINPUT89), .A3(new_n524_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n517_), .A2(new_n524_), .B1(KEYINPUT89), .B2(new_n502_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n451_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n502_), .A2(KEYINPUT89), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n522_), .A2(new_n523_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n522_), .A2(new_n523_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n517_), .A2(new_n524_), .A3(KEYINPUT89), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n449_), .A3(new_n450_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G8gat), .B(G36gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT18), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G64gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n217_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n406_), .A2(new_n401_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n396_), .A2(KEYINPUT90), .A3(new_n397_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542_));
  AND2_X1   g341(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n546_), .B2(new_n399_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n395_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n547_), .B2(new_n395_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n415_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n539_), .B1(new_n551_), .B2(new_n471_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT19), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n471_), .A2(new_n420_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n539_), .B1(new_n471_), .B2(new_n420_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n415_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n547_), .B2(new_n395_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n561_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n554_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n538_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n555_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n558_), .B(new_n555_), .C1(new_n551_), .C2(new_n471_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n538_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n550_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n547_), .A2(new_n548_), .A3(new_n395_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n560_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n471_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n556_), .B(KEYINPUT20), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n554_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n538_), .A3(new_n566_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n538_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT93), .B(KEYINPUT27), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n569_), .A2(KEYINPUT27), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n446_), .A2(new_n495_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT4), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n510_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n446_), .A2(new_n495_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(KEYINPUT4), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G225gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G1gat), .B(G29gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(G85gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT0), .ZN(new_n596_));
  INV_X1    g395(.A(G57gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n592_), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n534_), .A2(new_n582_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(KEYINPUT33), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n591_), .A2(new_n606_), .A3(new_n598_), .A4(new_n592_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n586_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n609_), .A2(new_n583_), .A3(KEYINPUT92), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT92), .B1(new_n609_), .B2(new_n583_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n590_), .A3(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n599_), .A3(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n608_), .A2(new_n576_), .A3(new_n578_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n557_), .A2(new_n563_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n538_), .A2(KEYINPUT32), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n575_), .A2(new_n566_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n618_), .B(new_n602_), .C1(new_n619_), .C2(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n525_), .A2(new_n526_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n451_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n604_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n387_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n355_), .A2(new_n361_), .A3(new_n343_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G8gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n308_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n362_), .A2(new_n633_), .A3(new_n365_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n310_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n630_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n308_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n310_), .A3(new_n639_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT75), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n641_), .B(KEYINPUT17), .C1(new_n644_), .C2(new_n630_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT76), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT17), .ZN(new_n647_));
  INV_X1    g446(.A(new_n630_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n637_), .A2(new_n640_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n647_), .B(new_n648_), .C1(new_n649_), .C2(KEYINPUT75), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n645_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n646_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n299_), .A2(new_n625_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n356_), .A3(new_n602_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT38), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n645_), .A2(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n294_), .A2(new_n296_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n625_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n356_), .B1(new_n659_), .B2(new_n602_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT94), .ZN(G1324gat));
  INV_X1    g461(.A(new_n582_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n343_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n654_), .B(new_n663_), .C1(new_n346_), .C2(new_n345_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT95), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g469(.A(new_n451_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n349_), .B1(new_n659_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT41), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n654_), .A2(new_n349_), .A3(new_n671_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(new_n622_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n350_), .B1(new_n659_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT42), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n350_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT96), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n654_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1327gat));
  NAND4_X1  g481(.A1(new_n653_), .A2(new_n337_), .A3(new_n385_), .A4(new_n341_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT97), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT37), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n658_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n294_), .A2(KEYINPUT37), .A3(new_n296_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n624_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n686_), .A2(new_n624_), .A3(new_n690_), .A4(new_n687_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n684_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(new_n684_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n690_), .B1(new_n299_), .B2(new_n624_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n691_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT98), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n692_), .A2(new_n700_), .A3(KEYINPUT44), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n602_), .B(new_n693_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT99), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(KEYINPUT98), .A3(new_n698_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n602_), .A4(new_n693_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(G29gat), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n703_), .A2(KEYINPUT100), .A3(G29gat), .A4(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n658_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n653_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n387_), .A3(new_n624_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT101), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n240_), .A3(new_n602_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT102), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n722_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1328gat));
  OR2_X1    g523(.A1(new_n582_), .A2(KEYINPUT103), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n582_), .A2(KEYINPUT103), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n241_), .A3(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT45), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n706_), .A2(new_n663_), .A3(new_n693_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n241_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1329gat));
  INV_X1    g533(.A(new_n718_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n243_), .B1(new_n735_), .B2(new_n451_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n706_), .A2(G43gat), .A3(new_n693_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n451_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n718_), .B2(new_n676_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n239_), .B(new_n622_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n693_), .ZN(G1331gat));
  AOI21_X1  g541(.A(new_n385_), .B1(new_n604_), .B2(new_n623_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n342_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n597_), .A3(new_n603_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n299_), .A2(new_n653_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n342_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT105), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(KEYINPUT105), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n743_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n602_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n746_), .B1(new_n753_), .B2(new_n597_), .ZN(G1332gat));
  OAI21_X1  g553(.A(G64gat), .B1(new_n745_), .B2(new_n727_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT106), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n758_), .A3(new_n728_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n761_), .A3(new_n671_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G71gat), .B1(new_n745_), .B2(new_n451_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT49), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1334gat));
  INV_X1    g564(.A(G78gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n752_), .A2(new_n766_), .A3(new_n676_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G78gat), .B1(new_n745_), .B2(new_n622_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT50), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1335gat));
  AND2_X1   g569(.A1(new_n744_), .A2(new_n716_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n602_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n342_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n715_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n386_), .B(new_n774_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT107), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n603_), .A2(new_n216_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n776_), .B2(new_n777_), .ZN(G1336gat));
  AOI21_X1  g577(.A(G92gat), .B1(new_n771_), .B2(new_n663_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n728_), .A2(G92gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT108), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT109), .ZN(G1337gat));
  AOI21_X1  g582(.A(new_n202_), .B1(new_n776_), .B2(new_n671_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n451_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n771_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n786_), .A2(KEYINPUT110), .A3(new_n787_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n786_), .A2(KEYINPUT111), .A3(new_n787_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT111), .B1(new_n786_), .B2(new_n787_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n790_), .A2(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(G1338gat));
  OAI21_X1  g593(.A(G106gat), .B1(new_n775_), .B2(new_n622_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT52), .B1(new_n795_), .B2(new_n796_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n797_), .B(new_n798_), .Z(new_n799_));
  NAND3_X1  g598(.A1(new_n771_), .A2(new_n207_), .A3(new_n676_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g601(.A1(new_n747_), .A2(new_n386_), .A3(new_n773_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n335_), .B2(KEYINPUT114), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n327_), .A2(new_n302_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n335_), .B2(KEYINPUT115), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n807_), .B(new_n808_), .C1(new_n806_), .C2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n339_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n339_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n329_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n375_), .B(KEYINPUT116), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n371_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n370_), .A2(new_n372_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n817_), .B(new_n381_), .C1(new_n371_), .C2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n384_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(KEYINPUT58), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n814_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n328_), .B(new_n820_), .C1(new_n822_), .C2(new_n812_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n299_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n385_), .A2(new_n328_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT113), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n822_), .B2(new_n812_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n820_), .B1(new_n336_), .B2(new_n329_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n827_), .B1(new_n832_), .B2(new_n714_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT57), .B(new_n658_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n826_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n805_), .B1(new_n835_), .B2(new_n657_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n663_), .A2(new_n603_), .A3(new_n533_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT117), .Z(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n385_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n835_), .A2(new_n657_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n842_), .B2(new_n805_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT59), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n835_), .A2(new_n653_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n845_), .B(new_n838_), .C1(new_n846_), .C2(new_n805_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT118), .B(G113gat), .Z(new_n849_));
  NOR2_X1   g648(.A1(new_n386_), .A2(new_n849_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT119), .Z(new_n851_));
  AOI21_X1  g650(.A(new_n841_), .B1(new_n848_), .B2(new_n851_), .ZN(G1340gat));
  OAI211_X1 g651(.A(new_n847_), .B(new_n342_), .C1(new_n840_), .C2(new_n845_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n844_), .A2(KEYINPUT120), .A3(new_n342_), .A4(new_n847_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(G120gat), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n438_), .B1(new_n773_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n840_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n438_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n840_), .B2(new_n715_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n645_), .A2(G127gat), .A3(new_n650_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n848_), .B2(new_n862_), .ZN(G1342gat));
  INV_X1    g662(.A(new_n299_), .ZN(new_n864_));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n847_), .B(new_n866_), .C1(new_n840_), .C2(new_n845_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n836_), .A2(new_n714_), .A3(new_n839_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT121), .B1(new_n868_), .B2(G134gat), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n865_), .C1(new_n843_), .C2(new_n714_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n869_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n867_), .A2(new_n869_), .A3(new_n871_), .A4(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1343gat));
  NOR4_X1   g675(.A1(new_n836_), .A2(new_n603_), .A3(new_n527_), .A4(new_n728_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n385_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n342_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n715_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n658_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n299_), .A2(G162gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT123), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n877_), .B2(new_n887_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n727_), .A2(new_n602_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n533_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n846_), .B2(new_n805_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n385_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n889_), .B1(new_n895_), .B2(G169gat), .ZN(new_n896_));
  AOI211_X1 g695(.A(KEYINPUT62), .B(new_n378_), .C1(new_n894_), .C2(new_n385_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT22), .B(G169gat), .Z(new_n898_));
  NOR2_X1   g697(.A1(new_n386_), .A2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT124), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n896_), .A2(new_n897_), .B1(new_n893_), .B2(new_n900_), .ZN(G1348gat));
  NOR3_X1   g700(.A1(new_n836_), .A2(new_n533_), .A3(new_n891_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(G176gat), .A3(new_n342_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n904_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n894_), .B2(new_n342_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1349gat));
  AOI21_X1  g707(.A(G183gat), .B1(new_n902_), .B2(new_n715_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n893_), .A2(new_n657_), .A3(new_n546_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n893_), .B2(new_n864_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n658_), .A2(new_n399_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n893_), .B2(new_n913_), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n836_), .A2(new_n527_), .A3(new_n891_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n385_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n342_), .A3(new_n458_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(new_n915_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G204gat), .B1(new_n920_), .B2(new_n773_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(G1353gat));
  NOR4_X1   g722(.A1(new_n836_), .A2(new_n657_), .A3(new_n527_), .A4(new_n891_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n928_), .A2(KEYINPUT127), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(KEYINPUT127), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n924_), .A2(new_n926_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1354gat));
  AOI21_X1  g731(.A(G218gat), .B1(new_n915_), .B2(new_n658_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n299_), .A2(G218gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n915_), .B2(new_n934_), .ZN(G1355gat));
endmodule


