//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT77), .ZN(new_n203_));
  OR3_X1    g002(.A1(new_n203_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n208_));
  OAI211_X1 g007(.A(KEYINPUT78), .B(new_n208_), .C1(new_n203_), .C2(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT22), .B(G169gat), .Z(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(G176gat), .C2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G197gat), .B(G204gat), .Z(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n203_), .A2(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  MUX2_X1   g026(.A(new_n226_), .B(KEYINPUT24), .S(new_n227_), .Z(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT26), .B(G190gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT91), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n225_), .B(new_n228_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n213_), .A2(new_n221_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n229_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n230_), .ZN(new_n235_));
  AND4_X1   g034(.A1(new_n209_), .A2(new_n204_), .A3(new_n228_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237_));
  INV_X1    g036(.A(G169gat), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT22), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT22), .B1(new_n237_), .B2(new_n238_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n211_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n225_), .B2(new_n207_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n220_), .B1(new_n236_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n245_), .A3(KEYINPUT20), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n244_), .A2(new_n236_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n221_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n213_), .A2(new_n232_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n252_), .B(KEYINPUT20), .C1(new_n253_), .C2(new_n221_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n254_), .B2(new_n249_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n249_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n246_), .A2(new_n249_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n260_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n265_), .A3(KEYINPUT27), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n263_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n260_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT93), .A3(new_n265_), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n268_), .A2(KEYINPUT93), .A3(new_n260_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT98), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT98), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n270_), .A2(new_n271_), .A3(new_n275_), .A4(new_n272_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n267_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G141gat), .B(G148gat), .Z(new_n278_));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(KEYINPUT83), .A3(G155gat), .A4(G162gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(KEYINPUT1), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT3), .Z(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT2), .Z(new_n289_));
  OAI22_X1  g088(.A1(new_n287_), .A2(new_n289_), .B1(G155gat), .B2(G162gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n279_), .B1(G155gat), .B2(G162gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n278_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n285_), .B1(new_n293_), .B2(new_n282_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G22gat), .B(G50gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n282_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n284_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n221_), .B1(new_n302_), .B2(KEYINPUT29), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n303_), .A2(KEYINPUT86), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT86), .B1(new_n303_), .B2(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(KEYINPUT85), .A3(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G78gat), .B(G106gat), .Z(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT87), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT88), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n300_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n307_), .A2(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(KEYINPUT89), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n307_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n300_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n316_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n318_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n321_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n320_), .A2(new_n325_), .B1(new_n328_), .B2(new_n300_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n251_), .B(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G113gat), .B(G120gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G134gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT82), .B(G127gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n331_), .B(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  XOR2_X1   g138(.A(G71gat), .B(G99gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT31), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n339_), .B(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n336_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n294_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(new_n335_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n335_), .A2(new_n347_), .ZN(new_n348_));
  OAI22_X1  g147(.A1(new_n346_), .A2(new_n347_), .B1(new_n294_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n350_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n353_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n343_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n277_), .A2(new_n329_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n320_), .A2(new_n325_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n328_), .A2(new_n300_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n359_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n270_), .A2(new_n271_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n354_), .B(new_n358_), .C1(KEYINPUT95), .C2(KEYINPUT33), .ZN(new_n371_));
  INV_X1    g170(.A(new_n335_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n345_), .B(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n358_), .B1(new_n373_), .B2(new_n351_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT96), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT96), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n375_), .B(new_n376_), .C1(new_n351_), .C2(new_n349_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n262_), .A2(new_n263_), .A3(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT97), .ZN(new_n381_));
  INV_X1    g180(.A(new_n379_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n380_), .A2(KEYINPUT97), .B1(new_n255_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n362_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n367_), .A2(new_n277_), .B1(new_n385_), .B2(new_n329_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n343_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n364_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT13), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT68), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT65), .B(KEYINPUT12), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G57gat), .A2(G64gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G57gat), .A2(G64gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT11), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G57gat), .ZN(new_n396_));
  INV_X1    g195(.A(G64gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(G78gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G71gat), .ZN(new_n402_));
  INV_X1    g201(.A(G71gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G78gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n398_), .A2(new_n392_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT11), .A3(new_n402_), .A4(new_n404_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT64), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(G99gat), .ZN(new_n415_));
  INV_X1    g214(.A(G106gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G99gat), .A2(G106gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n417_), .A2(new_n420_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT8), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT8), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n429_), .A3(new_n426_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT10), .B(G99gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n416_), .ZN(new_n432_));
  AND3_X1   g231(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n424_), .A2(KEYINPUT9), .A3(new_n425_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n425_), .A2(KEYINPUT9), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n428_), .A2(new_n430_), .B1(new_n432_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n391_), .B1(new_n413_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G230gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n413_), .B2(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n432_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n430_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n429_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT12), .A3(new_n408_), .A4(new_n406_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n440_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n440_), .A2(new_n443_), .A3(KEYINPUT66), .A4(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n413_), .A2(new_n439_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n442_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT5), .B(G176gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G204gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G120gat), .B(G148gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(KEYINPUT67), .A3(new_n465_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n390_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n389_), .A2(KEYINPUT68), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G8gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n483_), .B(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G229gat), .A3(G233gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n483_), .A2(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500_));
  INV_X1    g299(.A(new_n494_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n491_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(KEYINPUT15), .A3(new_n494_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n483_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n499_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n497_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n497_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n474_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n388_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n439_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n495_), .A2(new_n447_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT34), .Z(new_n527_));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(KEYINPUT72), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n520_), .A2(new_n523_), .A3(KEYINPUT71), .ZN(new_n532_));
  INV_X1    g331(.A(new_n529_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n528_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n529_), .B2(KEYINPUT71), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n527_), .A2(new_n522_), .A3(new_n528_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n521_), .A2(new_n524_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n530_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G190gat), .B(G218gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n544_), .B(KEYINPUT37), .C1(new_n546_), .C2(new_n539_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n539_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n539_), .A2(new_n546_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n547_), .B1(new_n552_), .B2(KEYINPUT37), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n483_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(new_n413_), .Z(new_n556_));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT16), .B(G183gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n555_), .B(new_n409_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n562_), .B(KEYINPUT76), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n553_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n519_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n476_), .A3(new_n362_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT38), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT100), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n518_), .B(KEYINPUT99), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n552_), .A2(new_n567_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n388_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n362_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n574_), .B(new_n579_), .C1(new_n572_), .C2(new_n571_), .ZN(G1324gat));
  INV_X1    g379(.A(new_n277_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(new_n477_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT39), .ZN(new_n583_));
  INV_X1    g382(.A(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n583_), .B1(new_n585_), .B2(G8gat), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT39), .B(new_n477_), .C1(new_n584_), .C2(new_n581_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT40), .Z(G1325gat));
  NOR2_X1   g388(.A1(new_n577_), .A2(new_n343_), .ZN(new_n590_));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT101), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n590_), .A2(KEYINPUT101), .A3(new_n591_), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n570_), .A2(new_n591_), .A3(new_n387_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(G1326gat));
  OAI21_X1  g398(.A(G22gat), .B1(new_n577_), .B2(new_n329_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT42), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n329_), .A2(G22gat), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n601_), .B1(new_n569_), .B2(new_n602_), .ZN(G1327gat));
  INV_X1    g402(.A(new_n552_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n567_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n519_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(G29gat), .B1(new_n608_), .B2(new_n362_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT89), .B1(new_n317_), .B2(new_n319_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n323_), .A2(new_n324_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n366_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n277_), .A2(new_n612_), .A3(new_n578_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n385_), .A2(new_n329_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n343_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(KEYINPUT103), .A3(new_n364_), .A4(new_n553_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n553_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n616_), .B2(new_n364_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n567_), .B(new_n617_), .C1(new_n619_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n575_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n387_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n277_), .A2(new_n329_), .A3(new_n363_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n625_), .B(new_n553_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n621_), .B1(new_n628_), .B2(new_n620_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n623_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT44), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(G29gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n622_), .B1(new_n388_), .B2(new_n553_), .ZN(new_n633_));
  NOR4_X1   g432(.A1(new_n626_), .A2(new_n625_), .A3(new_n627_), .A4(new_n618_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n605_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n628_), .A2(new_n620_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n575_), .A4(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n623_), .A2(new_n629_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n641_), .A2(KEYINPUT104), .A3(KEYINPUT44), .A4(new_n575_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n578_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n609_), .B1(new_n632_), .B2(new_n643_), .ZN(G1328gat));
  INV_X1    g443(.A(G36gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n608_), .A2(new_n645_), .A3(new_n581_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT45), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n581_), .B1(new_n630_), .B2(KEYINPUT44), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n649_), .B2(new_n645_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT46), .B(new_n647_), .C1(new_n649_), .C2(new_n645_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND2_X1  g453(.A1(new_n640_), .A2(new_n642_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n655_), .A2(G43gat), .A3(new_n387_), .A4(new_n631_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT105), .B(G43gat), .Z(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n607_), .B2(new_n343_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT106), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT47), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1330gat));
  INV_X1    g463(.A(G50gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n608_), .A2(new_n665_), .A3(new_n612_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n329_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n667_), .B(new_n665_), .C1(new_n668_), .C2(new_n631_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n655_), .A2(new_n612_), .A3(new_n631_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n670_), .B2(G50gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n669_), .B2(new_n671_), .ZN(G1331gat));
  NAND2_X1  g471(.A1(new_n474_), .A2(new_n517_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n616_), .B2(new_n364_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n576_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(new_n396_), .A3(new_n578_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n568_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n362_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n396_), .B2(new_n679_), .ZN(G1332gat));
  OAI21_X1  g479(.A(G64gat), .B1(new_n675_), .B2(new_n277_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT108), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT48), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n397_), .A3(new_n581_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(G1333gat));
  OAI21_X1  g486(.A(G71gat), .B1(new_n675_), .B2(new_n343_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT49), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n678_), .A2(new_n403_), .A3(new_n387_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1334gat));
  OAI21_X1  g490(.A(G78gat), .B1(new_n675_), .B2(new_n329_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT50), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n401_), .A3(new_n612_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1335gat));
  NAND2_X1  g494(.A1(new_n674_), .A2(new_n606_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n362_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n623_), .A2(new_n629_), .A3(new_n673_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n578_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n698_), .B1(new_n701_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g501(.A(G92gat), .B1(new_n697_), .B2(new_n581_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n581_), .A2(G92gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n699_), .B2(new_n704_), .ZN(G1337gat));
  OAI21_X1  g504(.A(G99gat), .B1(new_n700_), .B2(new_n343_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n431_), .A3(new_n387_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g508(.A(new_n416_), .B1(new_n699_), .B2(new_n612_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT52), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT52), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n696_), .A2(G106gat), .A3(new_n329_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT109), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n712_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n711_), .A2(new_n717_), .A3(new_n712_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  NAND2_X1  g518(.A1(new_n516_), .A2(new_n465_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n440_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n440_), .A2(new_n448_), .A3(KEYINPUT111), .A4(new_n455_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n442_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n428_), .A2(new_n430_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n409_), .B1(new_n728_), .B2(new_n444_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n454_), .A2(new_n391_), .B1(new_n729_), .B2(KEYINPUT12), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT66), .B1(new_n730_), .B2(new_n443_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n452_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n449_), .A2(new_n727_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(KEYINPUT56), .A3(new_n462_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT113), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n736_), .A2(new_n739_), .A3(KEYINPUT56), .A4(new_n462_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n462_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(KEYINPUT56), .C1(new_n736_), .C2(new_n462_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n720_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n496_), .A2(new_n499_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n498_), .A2(new_n507_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n749_), .B(new_n512_), .C1(new_n750_), .C2(new_n499_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(new_n515_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n468_), .A2(new_n752_), .A3(new_n469_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT57), .B(new_n604_), .C1(new_n748_), .C2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT115), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT55), .B1(new_n451_), .B2(new_n452_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n441_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n464_), .B1(new_n759_), .B2(new_n735_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n745_), .B1(new_n760_), .B2(KEYINPUT56), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n757_), .A2(new_n758_), .A3(new_n734_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT112), .B(new_n743_), .C1(new_n762_), .C2(new_n464_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n761_), .A2(new_n738_), .A3(new_n740_), .A4(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n720_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n552_), .B1(new_n766_), .B2(new_n753_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT57), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n756_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n737_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n736_), .B2(new_n462_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n465_), .B(new_n752_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n737_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT58), .A3(new_n465_), .A4(new_n752_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n778_), .A3(new_n553_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n754_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n552_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n567_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT119), .ZN(new_n785_));
  INV_X1    g584(.A(new_n474_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n517_), .A3(new_n568_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n783_), .A2(new_n790_), .A3(new_n567_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n277_), .A2(new_n362_), .A3(new_n329_), .A4(new_n387_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT118), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n768_), .B1(new_n767_), .B2(KEYINPUT57), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n781_), .A2(KEYINPUT115), .A3(new_n780_), .A4(new_n552_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n779_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n775_), .A2(new_n778_), .A3(new_n553_), .A4(KEYINPUT114), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n782_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n798_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n803_), .A2(new_n782_), .A3(new_n804_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n770_), .A2(new_n807_), .A3(KEYINPUT116), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n567_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n789_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(new_n789_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n795_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n797_), .B1(new_n814_), .B2(KEYINPUT59), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(G113gat), .A3(new_n516_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n814_), .B2(new_n517_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1340gat));
  AND2_X1   g618(.A1(new_n813_), .A2(new_n795_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n474_), .B(new_n796_), .C1(new_n820_), .C2(new_n793_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n786_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n820_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n814_), .B2(new_n567_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n827_), .C1(new_n814_), .C2(new_n567_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n567_), .A2(new_n827_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n796_), .B(new_n832_), .C1(new_n820_), .C2(new_n793_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .ZN(G1342gat));
  AOI21_X1  g633(.A(G134gat), .B1(new_n820_), .B2(new_n552_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT121), .B(G134gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n618_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n815_), .B2(new_n837_), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n809_), .A2(new_n789_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n809_), .A2(new_n810_), .A3(new_n789_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n581_), .A2(new_n578_), .A3(new_n329_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n840_), .A2(new_n343_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n517_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n786_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g646(.A1(new_n843_), .A2(new_n567_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  NOR3_X1   g649(.A1(new_n811_), .A2(new_n812_), .A3(new_n387_), .ZN(new_n851_));
  INV_X1    g650(.A(G162gat), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n552_), .A4(new_n842_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G162gat), .B1(new_n843_), .B2(new_n618_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1347gat));
  NAND2_X1  g657(.A1(new_n581_), .A2(new_n363_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n517_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT123), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(KEYINPUT123), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n792_), .A2(new_n329_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n863_), .A2(new_n864_), .A3(G169gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(G169gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n792_), .A2(new_n329_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n859_), .A2(new_n517_), .A3(new_n212_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n865_), .A2(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n859_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n792_), .A2(new_n474_), .A3(new_n329_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n240_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n813_), .B2(new_n329_), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT125), .A4(new_n612_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n474_), .A2(G176gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n873_), .B1(new_n879_), .B2(new_n870_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n867_), .A2(new_n859_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n881_), .A2(new_n231_), .A3(new_n605_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n605_), .B(new_n870_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n205_), .ZN(G1350gat));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n234_), .A3(new_n552_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n553_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(G190gat), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT126), .B(new_n206_), .C1(new_n881_), .C2(new_n553_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1351gat));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n277_), .A2(new_n329_), .A3(new_n362_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n813_), .A2(new_n891_), .A3(new_n343_), .A4(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n840_), .A2(new_n343_), .A3(new_n841_), .A4(new_n892_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT127), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G197gat), .B1(new_n896_), .B2(new_n516_), .ZN(new_n897_));
  INV_X1    g696(.A(G197gat), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n898_), .B(new_n517_), .C1(new_n893_), .C2(new_n895_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1352gat));
  AOI21_X1  g699(.A(G204gat), .B1(new_n896_), .B2(new_n474_), .ZN(new_n901_));
  INV_X1    g700(.A(G204gat), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n902_), .B(new_n786_), .C1(new_n893_), .C2(new_n895_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1353gat));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n567_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n896_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n907_), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n905_), .B(new_n909_), .C1(new_n893_), .C2(new_n895_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1354gat));
  AOI21_X1  g710(.A(G218gat), .B1(new_n896_), .B2(new_n552_), .ZN(new_n912_));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n913_), .B(new_n618_), .C1(new_n893_), .C2(new_n895_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1355gat));
endmodule


