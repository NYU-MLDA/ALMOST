//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n210_), .B(new_n211_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n213_), .B(new_n214_), .C1(G99gat), .C2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT65), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n209_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  AND2_X1   g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n219_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n225_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n212_), .A2(new_n215_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT8), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT64), .B(G92gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(G85gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n211_), .A3(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n234_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n217_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT65), .B1(new_n204_), .B2(new_n206_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n228_), .A2(new_n231_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G29gat), .B(G36gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G43gat), .B(G50gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n244_), .A2(new_n245_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n245_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n202_), .B1(new_n243_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT34), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n252_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n243_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n249_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n246_), .A2(new_n247_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n248_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n216_), .A2(new_n207_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n225_), .A3(new_n222_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n266_), .A2(KEYINPUT8), .B1(new_n218_), .B2(new_n227_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n234_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n268_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n264_), .B(KEYINPUT72), .C1(new_n267_), .C2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n255_), .A2(new_n260_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n256_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT70), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(new_n276_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n278_), .A2(KEYINPUT70), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT75), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n277_), .A2(new_n279_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n243_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n264_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n271_), .A2(new_n280_), .B1(new_n288_), .B2(new_n260_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G190gat), .B(G218gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT73), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G134gat), .B(G162gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT36), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(KEYINPUT36), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n289_), .A2(KEYINPUT74), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n289_), .B2(KEYINPUT74), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  NOR2_X1   g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  MUX2_X1   g102(.A(new_n302_), .B(new_n303_), .S(KEYINPUT86), .Z(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT31), .Z(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT23), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT22), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(KEYINPUT22), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n319_), .B(new_n322_), .C1(new_n323_), .C2(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n318_), .A2(KEYINPUT24), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n328_), .B(new_n331_), .C1(new_n329_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n311_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n313_), .A2(KEYINPUT82), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n313_), .A2(KEYINPUT82), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n325_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G99gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(G71gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n339_), .B(new_n210_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n308_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n347_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n307_), .A3(new_n350_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(G141gat), .ZN(new_n366_));
  INV_X1    g165(.A(G148gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT3), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n365_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT87), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n371_), .A2(KEYINPUT89), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT89), .B1(new_n371_), .B2(new_n377_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n364_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n361_), .A2(KEYINPUT1), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n363_), .B1(new_n362_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n373_), .B(new_n375_), .C1(G141gat), .C2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n360_), .B1(new_n380_), .B2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G197gat), .B(G204gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(KEYINPUT21), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n359_), .B1(new_n390_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n387_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n368_), .A2(new_n370_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n365_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n377_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n371_), .A2(KEYINPUT89), .A3(new_n377_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n402_), .B1(new_n409_), .B2(new_n364_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n399_), .B(new_n358_), .C1(new_n410_), .C2(new_n360_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT91), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n401_), .B2(new_n411_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(KEYINPUT92), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  AOI211_X1 g216(.A(new_n417_), .B(new_n413_), .C1(new_n401_), .C2(new_n411_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G22gat), .B(G50gat), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n380_), .A2(new_n360_), .A3(new_n389_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT28), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT28), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n380_), .A2(new_n425_), .A3(new_n360_), .A4(new_n389_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n410_), .B2(new_n360_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n426_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT90), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n420_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT93), .B1(new_n419_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n413_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n390_), .A2(new_n400_), .A3(new_n359_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n364_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT29), .B1(new_n440_), .B2(new_n402_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n358_), .B1(new_n441_), .B2(new_n399_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n437_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n417_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n415_), .A2(KEYINPUT92), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n414_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n427_), .A2(new_n428_), .A3(new_n421_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n420_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT93), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n436_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n443_), .A2(new_n414_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n434_), .B2(new_n429_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT94), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT94), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n457_), .B(new_n454_), .C1(new_n436_), .C2(new_n451_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n357_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n419_), .A2(KEYINPUT93), .A3(new_n435_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n450_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n455_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n457_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(KEYINPUT94), .A3(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n353_), .A2(new_n356_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n321_), .A2(KEYINPUT22), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n323_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n318_), .B1(new_n473_), .B2(G176gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n337_), .A2(new_n475_), .A3(new_n315_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n337_), .B2(new_n315_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n314_), .A2(new_n331_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT97), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n329_), .B1(new_n332_), .B2(KEYINPUT96), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(KEYINPUT96), .B2(new_n332_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n328_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n399_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  INV_X1    g284(.A(new_n338_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n400_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n470_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT20), .B1(new_n400_), .B2(new_n486_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n478_), .A2(new_n483_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n400_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n488_), .A2(new_n489_), .B1(new_n493_), .B2(new_n470_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G8gat), .B(G36gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n490_), .A2(new_n494_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n467_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n490_), .A2(new_n494_), .A3(new_n500_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(new_n470_), .A3(new_n487_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n493_), .B2(new_n470_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n506_), .A2(KEYINPUT103), .A3(new_n499_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT103), .B1(new_n506_), .B2(new_n499_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n504_), .B(KEYINPUT27), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n380_), .A2(new_n389_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n304_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n302_), .B2(new_n511_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT4), .B1(new_n304_), .B2(new_n511_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n513_), .B2(KEYINPUT4), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G225gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  MUX2_X1   g316(.A(new_n513_), .B(new_n515_), .S(new_n517_), .Z(new_n518_));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G85gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n513_), .A2(new_n516_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n510_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n459_), .A2(new_n466_), .A3(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n456_), .A2(new_n458_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n490_), .A2(new_n494_), .A3(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n506_), .A2(KEYINPUT32), .A3(new_n500_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n526_), .A2(new_n527_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT33), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n513_), .A2(new_n516_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n527_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT102), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(KEYINPUT102), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n538_), .A2(new_n541_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n501_), .A2(new_n502_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n536_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n532_), .A2(new_n547_), .A3(new_n465_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n299_), .B1(new_n531_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(G64gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G57gat), .ZN(new_n551_));
  INV_X1    g350(.A(G57gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G64gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT11), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n553_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT69), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT11), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n342_), .A2(KEYINPUT68), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G71gat), .ZN(new_n565_));
  INV_X1    g364(.A(G78gat), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n558_), .A2(new_n562_), .A3(new_n569_), .ZN(new_n570_));
  OAI221_X1 g369(.A(KEYINPUT11), .B1(new_n567_), .B2(new_n568_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n570_), .B(new_n571_), .C1(new_n267_), .C2(new_n269_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n243_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n574_), .A3(KEYINPUT12), .ZN(new_n575_));
  OR3_X1    g374(.A1(new_n243_), .A2(new_n573_), .A3(KEYINPUT12), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n578_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n589_), .B2(new_n580_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT13), .B1(new_n587_), .B2(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n573_), .B(new_n597_), .Z(new_n598_));
  XNOR2_X1  g397(.A(G1gat), .B(G8gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT78), .B(G15gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G22gat), .ZN(new_n602_));
  INV_X1    g401(.A(G22gat), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(G15gat), .ZN(new_n605_));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT78), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT14), .ZN(new_n610_));
  INV_X1    g409(.A(G1gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT79), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT79), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G1gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n610_), .B1(new_n615_), .B2(G8gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n600_), .B1(new_n609_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT79), .B(G1gat), .ZN(new_n618_));
  INV_X1    g417(.A(G8gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT14), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(new_n602_), .A3(new_n608_), .A4(new_n599_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n598_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n623_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n623_), .A2(new_n629_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n617_), .A2(new_n262_), .A3(new_n621_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT81), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n622_), .B2(new_n259_), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT81), .B(new_n262_), .C1(new_n617_), .C2(new_n621_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n635_), .B(new_n637_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n254_), .A2(new_n622_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n622_), .A2(new_n259_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT81), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n622_), .A2(new_n638_), .A3(new_n259_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n646_), .B2(new_n637_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G169gat), .B(G197gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n648_), .B(new_n649_), .Z(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n641_), .B(new_n652_), .C1(new_n646_), .C2(new_n637_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n596_), .A2(new_n634_), .A3(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n549_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n529_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n531_), .A2(new_n548_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT104), .B1(new_n661_), .B2(new_n654_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n663_), .B(new_n655_), .C1(new_n531_), .C2(new_n548_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT37), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT76), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT77), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n289_), .A2(new_n294_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n271_), .A2(new_n280_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n288_), .A2(new_n260_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(KEYINPUT74), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n296_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n289_), .A2(KEYINPUT74), .A3(new_n296_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n670_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n666_), .A2(KEYINPUT76), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n669_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n299_), .A2(new_n680_), .A3(new_n668_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n633_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n596_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n529_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n529_), .A2(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n615_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n665_), .A2(new_n684_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n692_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n660_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT107), .ZN(G1324gat));
  AND2_X1   g495(.A1(new_n665_), .A2(new_n684_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n619_), .A3(new_n510_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n510_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G8gat), .B1(new_n658_), .B2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT39), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT39), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1325gat));
  AOI21_X1  g504(.A(new_n606_), .B1(new_n657_), .B2(new_n357_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT41), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n697_), .A2(new_n606_), .A3(new_n357_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1326gat));
  INV_X1    g508(.A(new_n532_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n603_), .B1(new_n657_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n697_), .A2(new_n603_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1327gat));
  NOR3_X1   g514(.A1(new_n596_), .A2(new_n633_), .A3(new_n655_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n682_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT43), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n661_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n682_), .B1(new_n531_), .B2(new_n548_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n716_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT44), .B(new_n716_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G29gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n689_), .A2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n596_), .A2(new_n677_), .A3(new_n633_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT110), .B(new_n731_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n529_), .A3(new_n735_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n728_), .A2(new_n730_), .B1(new_n736_), .B2(new_n729_), .ZN(G1328gat));
  NOR2_X1   g536(.A1(new_n699_), .A2(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n735_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT45), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n734_), .A2(new_n741_), .A3(new_n735_), .A4(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n510_), .A3(new_n727_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G36gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(KEYINPUT46), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1329gat));
  NAND3_X1  g549(.A1(new_n728_), .A2(G43gat), .A3(new_n357_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n734_), .A2(new_n357_), .A3(new_n735_), .ZN(new_n752_));
  INV_X1    g551(.A(G43gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n757_), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1330gat));
  INV_X1    g558(.A(G50gat), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n532_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n734_), .A2(new_n710_), .A3(new_n735_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n728_), .A2(new_n761_), .B1(new_n762_), .B2(new_n760_), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n683_), .A2(new_n595_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n654_), .B1(new_n531_), .B2(new_n548_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n689_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G57gat), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  AND4_X1   g568(.A1(new_n549_), .A2(new_n633_), .A3(new_n655_), .A4(new_n596_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT112), .B(G57gat), .Z(new_n771_));
  NOR2_X1   g570(.A1(new_n659_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n769_), .B1(new_n770_), .B2(new_n772_), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n550_), .B1(new_n770_), .B2(new_n510_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT48), .Z(new_n775_));
  NAND3_X1  g574(.A1(new_n767_), .A2(new_n550_), .A3(new_n510_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1333gat));
  AOI21_X1  g576(.A(new_n342_), .B1(new_n770_), .B2(new_n357_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT49), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n767_), .A2(new_n342_), .A3(new_n357_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1334gat));
  AOI21_X1  g580(.A(new_n566_), .B1(new_n770_), .B2(new_n710_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT50), .Z(new_n783_));
  NAND3_X1  g582(.A1(new_n767_), .A2(new_n566_), .A3(new_n710_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1335gat));
  AND4_X1   g584(.A1(new_n299_), .A2(new_n766_), .A3(new_n634_), .A4(new_n596_), .ZN(new_n786_));
  INV_X1    g585(.A(G85gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n768_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n596_), .A2(new_n634_), .A3(new_n655_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n721_), .A2(new_n722_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n721_), .A2(new_n719_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT113), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n789_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n529_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n796_), .B2(new_n787_), .ZN(G1336gat));
  AOI21_X1  g596(.A(G92gat), .B1(new_n786_), .B2(new_n510_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n510_), .A2(new_n232_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n795_), .B2(new_n799_), .ZN(G1337gat));
  NAND4_X1  g599(.A1(new_n786_), .A2(new_n236_), .A3(new_n237_), .A4(new_n357_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n795_), .A2(new_n357_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n210_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT51), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n801_), .C1(new_n802_), .C2(new_n210_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n532_), .A2(new_n789_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G106gat), .B1(new_n808_), .B2(KEYINPUT114), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n811_), .A2(KEYINPUT114), .A3(new_n808_), .A4(G106gat), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n532_), .A2(G106gat), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n814_), .A2(new_n815_), .B1(new_n786_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n817_), .B(new_n819_), .ZN(G1339gat));
  NAND4_X1  g619(.A1(new_n682_), .A2(new_n633_), .A3(new_n655_), .A4(new_n595_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT54), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n575_), .A2(new_n576_), .A3(new_n588_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n823_), .A2(new_n589_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n577_), .A2(new_n824_), .A3(new_n578_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n585_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n825_), .A2(new_n827_), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n589_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n653_), .B2(new_n651_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n575_), .A2(new_n576_), .A3(new_n588_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n579_), .A2(KEYINPUT55), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n586_), .B1(new_n589_), .B2(new_n824_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n828_), .A2(new_n830_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n650_), .B1(new_n839_), .B2(new_n636_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n646_), .A2(new_n637_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n647_), .A2(new_n650_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n586_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(KEYINPUT118), .C1(new_n843_), .C2(new_n829_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n591_), .B2(new_n842_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n828_), .A2(new_n830_), .A3(KEYINPUT117), .A4(new_n835_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n677_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT57), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n852_), .A3(new_n677_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n827_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n587_), .A3(new_n842_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n825_), .A2(new_n827_), .A3(KEYINPUT56), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(KEYINPUT58), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n682_), .B1(KEYINPUT58), .B2(new_n857_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n851_), .A2(new_n853_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n822_), .B1(new_n860_), .B2(new_n633_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n689_), .A2(new_n510_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n532_), .A3(new_n357_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n634_), .B1(new_n860_), .B2(KEYINPUT120), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n822_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(new_n865_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n871_), .B2(new_n862_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872_), .B2(new_n655_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n874_), .A3(new_n654_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1340gat));
  OAI21_X1  g675(.A(G120gat), .B1(new_n872_), .B2(new_n595_), .ZN(new_n877_));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n595_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n871_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n878_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n872_), .B2(new_n634_), .ZN(new_n882_));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n883_), .A3(new_n633_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1342gat));
  OAI21_X1  g684(.A(G134gat), .B1(new_n872_), .B2(new_n682_), .ZN(new_n886_));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n871_), .A2(new_n887_), .A3(new_n299_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n532_), .A2(new_n357_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n870_), .A2(new_n863_), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n655_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n366_), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n595_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n367_), .ZN(G1345gat));
  INV_X1    g694(.A(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n633_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  OR3_X1    g698(.A1(new_n891_), .A2(G162gat), .A3(new_n677_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n891_), .B2(new_n682_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n821_), .B(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n859_), .A2(new_n858_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n849_), .A2(new_n852_), .A3(new_n677_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n852_), .B1(new_n849_), .B2(new_n677_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n908_), .B2(new_n634_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n688_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n357_), .B1(new_n910_), .B2(new_n686_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT121), .B1(new_n911_), .B2(new_n699_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n689_), .A2(new_n913_), .A3(new_n357_), .A4(new_n510_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n710_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n909_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n321_), .B1(new_n917_), .B2(new_n654_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT62), .Z(new_n919_));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n909_), .B2(new_n916_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n851_), .A2(new_n853_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n633_), .B1(new_n922_), .B2(new_n905_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT122), .B(new_n915_), .C1(new_n923_), .C2(new_n904_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n472_), .A3(new_n654_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n919_), .A2(new_n926_), .ZN(G1348gat));
  NAND2_X1  g726(.A1(new_n912_), .A2(new_n914_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n595_), .A2(new_n319_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n870_), .A2(new_n532_), .A3(new_n928_), .A4(new_n929_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n909_), .A2(new_n916_), .A3(new_n920_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT122), .B1(new_n861_), .B2(new_n915_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n596_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n933_), .B2(new_n319_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n595_), .B1(new_n921_), .B2(new_n924_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n935_), .A2(new_n936_), .A3(G176gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n930_), .B1(new_n934_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT124), .B(new_n930_), .C1(new_n934_), .C2(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1349gat));
  NAND4_X1  g741(.A1(new_n870_), .A2(new_n532_), .A3(new_n633_), .A4(new_n928_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n634_), .A2(new_n326_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n943_), .A2(new_n309_), .B1(new_n925_), .B2(new_n944_), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n925_), .A2(new_n299_), .A3(new_n327_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n682_), .B1(new_n921_), .B2(new_n924_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n310_), .ZN(G1351gat));
  NOR2_X1   g747(.A1(new_n699_), .A2(new_n529_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n870_), .A2(new_n890_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n654_), .ZN(new_n951_));
  INV_X1    g750(.A(G197gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(KEYINPUT125), .B2(new_n952_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT125), .B(G197gat), .Z(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n951_), .B2(new_n954_), .ZN(G1352gat));
  AOI21_X1  g754(.A(new_n595_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n950_), .A2(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n957_), .B(new_n958_), .Z(G1353gat));
  NAND2_X1  g758(.A1(new_n950_), .A2(new_n633_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  AND2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n960_), .B2(new_n961_), .ZN(G1354gat));
  NOR2_X1   g763(.A1(new_n677_), .A2(G218gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n950_), .A2(new_n965_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n950_), .A2(new_n717_), .ZN(new_n967_));
  INV_X1    g766(.A(G218gat), .ZN(new_n968_));
  OAI211_X1 g767(.A(KEYINPUT127), .B(new_n966_), .C1(new_n967_), .C2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970_));
  INV_X1    g769(.A(new_n966_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n968_), .B1(new_n950_), .B2(new_n717_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n970_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n969_), .A2(new_n973_), .ZN(G1355gat));
endmodule


