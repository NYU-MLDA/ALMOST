//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n205_), .B2(KEYINPUT1), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(KEYINPUT1), .B2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT83), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n211_), .B(KEYINPUT3), .Z(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n209_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT85), .Z(new_n219_));
  AND2_X1   g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT86), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n213_), .B(new_n214_), .C1(new_n220_), .C2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n221_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n219_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n227_), .A2(new_n228_), .B1(new_n207_), .B2(new_n212_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n224_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n214_), .A3(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G22gat), .B(G50gat), .Z(new_n232_));
  AND3_X1   g031(.A1(new_n225_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G78gat), .B(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT92), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n233_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT88), .B(G197gat), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G204gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT21), .B1(new_n241_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G211gat), .B(G218gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT90), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G197gat), .A2(G204gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(new_n239_), .B2(G204gat), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n246_), .B(new_n248_), .C1(KEYINPUT21), .C2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n229_), .B2(new_n214_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n254_), .B2(KEYINPUT91), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  OAI221_X1 g057(.A(new_n254_), .B1(KEYINPUT91), .B2(new_n256_), .C1(new_n229_), .C2(new_n214_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n236_), .A3(new_n235_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n235_), .A2(new_n236_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n238_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n235_), .A2(KEYINPUT93), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n258_), .A2(new_n259_), .A3(KEYINPUT93), .A4(new_n235_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n266_), .B(new_n267_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(KEYINPUT23), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT23), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(KEYINPUT80), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(KEYINPUT80), .B2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(G183gat), .B2(G190gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n279_), .A2(KEYINPUT78), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(KEYINPUT78), .ZN(new_n281_));
  OAI21_X1  g080(.A(G190gat), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT25), .B(G183gat), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n279_), .A2(KEYINPUT77), .A3(G190gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT77), .B1(new_n279_), .B2(G190gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT79), .B1(new_n270_), .B2(KEYINPUT23), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(new_n272_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  NOR3_X1   g089(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n278_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT81), .B(G15gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n294_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT82), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n298_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305_));
  INV_X1    g104(.A(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT30), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n304_), .B(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n213_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n302_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n229_), .A2(new_n303_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT4), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT96), .Z(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT97), .B(KEYINPUT4), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n314_), .B(new_n316_), .C1(new_n312_), .C2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n312_), .A2(new_n313_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n319_), .A2(new_n326_), .A3(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n310_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n254_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n288_), .B1(G183gat), .B2(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n277_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT26), .B(G190gat), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n283_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n274_), .A2(new_n292_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n254_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n254_), .A2(new_n344_), .A3(KEYINPUT94), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n337_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n254_), .A2(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n294_), .A2(new_n254_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n354_), .A2(KEYINPUT20), .A3(new_n352_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n336_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n335_), .B(new_n356_), .C1(new_n349_), .C2(new_n352_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n353_), .A2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(KEYINPUT95), .A3(new_n335_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n349_), .A2(new_n352_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n354_), .A2(KEYINPUT20), .A3(new_n355_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n351_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n335_), .B(KEYINPUT98), .Z(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT27), .B(new_n360_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  AND4_X1   g170(.A1(new_n269_), .A2(new_n331_), .A3(new_n365_), .A4(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n269_), .A2(new_n330_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n363_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n312_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n327_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n312_), .A2(new_n318_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n320_), .B2(KEYINPUT4), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n379_), .B2(new_n315_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n329_), .A2(KEYINPUT33), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n319_), .A2(new_n382_), .A3(new_n321_), .A4(new_n326_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n362_), .B2(new_n385_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n375_), .A2(new_n384_), .B1(new_n330_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n269_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n374_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n372_), .B1(new_n390_), .B2(new_n310_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT10), .B(G99gat), .Z(new_n392_));
  INV_X1    g191(.A(G106gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G85gat), .B(G92gat), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT9), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT6), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G99gat), .A3(G106gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G85gat), .ZN(new_n402_));
  INV_X1    g201(.A(G92gat), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT9), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n394_), .A2(new_n396_), .A3(new_n401_), .A4(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT8), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(G99gat), .B2(G106gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n397_), .A2(KEYINPUT6), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT66), .ZN(new_n411_));
  INV_X1    g210(.A(G99gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n393_), .A3(KEYINPUT65), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT7), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n412_), .A3(new_n393_), .A4(KEYINPUT65), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n410_), .A2(new_n411_), .A3(new_n414_), .A4(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n406_), .B1(new_n417_), .B2(new_n395_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n401_), .A3(new_n416_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n406_), .A3(new_n395_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT69), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n424_), .B(new_n405_), .C1(new_n418_), .C2(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT12), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G57gat), .B(G64gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n430_), .A2(new_n431_), .A3(G78gat), .ZN(new_n432_));
  INV_X1    g231(.A(G64gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G57gat), .ZN(new_n434_));
  INV_X1    g233(.A(G57gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G64gat), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT11), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(G78gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n429_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n441_));
  INV_X1    g240(.A(G78gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n439_), .C1(KEYINPUT11), .C2(new_n427_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(KEYINPUT68), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n428_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(KEYINPUT68), .ZN(new_n448_));
  INV_X1    g247(.A(new_n437_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n429_), .A3(new_n439_), .A4(new_n444_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n428_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n426_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n423_), .A2(new_n425_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G230gat), .A2(G233gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT64), .Z(new_n456_));
  INV_X1    g255(.A(new_n405_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n417_), .A2(new_n395_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT8), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n459_), .B2(new_n420_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n451_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n426_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n460_), .A2(new_n463_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n454_), .B(new_n456_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n456_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n447_), .A2(new_n452_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(new_n422_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G120gat), .B(G148gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT5), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G176gat), .B(G204gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n475_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n466_), .A2(new_n470_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(KEYINPUT13), .A3(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G29gat), .B(G36gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT70), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n485_), .A2(KEYINPUT70), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(KEYINPUT70), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496_));
  INV_X1    g295(.A(G1gat), .ZN(new_n497_));
  INV_X1    g296(.A(G8gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G1gat), .B(G8gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(KEYINPUT15), .A3(new_n492_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n495_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n492_), .B2(new_n489_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT75), .ZN(new_n509_));
  INV_X1    g308(.A(new_n505_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n502_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n493_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(new_n506_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n504_), .A2(new_n514_), .A3(new_n505_), .A4(new_n507_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G113gat), .B(G141gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT76), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n509_), .A2(new_n513_), .A3(new_n515_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n484_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n391_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n502_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n468_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT16), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n529_), .A2(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(KEYINPUT17), .A3(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n489_), .A2(KEYINPUT15), .A3(new_n492_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT15), .B1(new_n489_), .B2(new_n492_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n423_), .A2(new_n546_), .A3(new_n425_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n460_), .A2(new_n493_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n548_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n547_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(KEYINPUT71), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n547_), .A2(new_n552_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n553_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n547_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n561_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n560_), .B(KEYINPUT36), .ZN(new_n571_));
  OAI221_X1 g370(.A(new_n569_), .B1(KEYINPUT72), .B2(new_n570_), .C1(new_n557_), .C2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT71), .B1(new_n557_), .B2(new_n561_), .ZN(new_n573_));
  AND4_X1   g372(.A1(KEYINPUT71), .A2(new_n564_), .A3(new_n565_), .A4(new_n561_), .ZN(new_n574_));
  OAI22_X1  g373(.A1(new_n573_), .A2(new_n574_), .B1(new_n557_), .B2(new_n571_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT72), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n543_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT74), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n526_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n330_), .A2(KEYINPUT100), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n330_), .A2(KEYINPUT100), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n580_), .A2(KEYINPUT101), .A3(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT101), .B1(new_n580_), .B2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT102), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .A4(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n589_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n557_), .A2(new_n571_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n568_), .B2(new_n562_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n391_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n525_), .A2(new_n543_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n330_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT103), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n594_), .A3(new_n602_), .ZN(G1324gat));
  NAND2_X1  g402(.A1(new_n365_), .A2(new_n371_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n526_), .A2(new_n498_), .A3(new_n604_), .A4(new_n579_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n599_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(G1325gat));
  OR3_X1    g411(.A1(new_n580_), .A2(G15gat), .A3(new_n310_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G15gat), .B1(new_n599_), .B2(new_n310_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT41), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1326gat));
  OAI21_X1  g419(.A(G22gat), .B1(new_n599_), .B2(new_n269_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT42), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n269_), .A2(G22gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n580_), .B2(new_n623_), .ZN(G1327gat));
  NOR2_X1   g423(.A1(new_n575_), .A2(new_n542_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n526_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G29gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n330_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n525_), .A2(KEYINPUT105), .A3(new_n542_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT105), .B1(new_n525_), .B2(new_n542_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n629_), .A2(new_n630_), .B1(KEYINPUT107), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n375_), .A2(new_n384_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n387_), .A2(new_n330_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n389_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n373_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n310_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n372_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n572_), .A2(new_n577_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n633_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n391_), .A2(KEYINPUT43), .A3(new_n641_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n632_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT107), .B1(new_n631_), .B2(KEYINPUT106), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n632_), .B(new_n648_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n583_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n628_), .B1(new_n650_), .B2(new_n627_), .ZN(G1328gat));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n604_), .B(KEYINPUT108), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n526_), .A2(new_n652_), .A3(new_n625_), .A4(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n606_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n652_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n656_), .B(new_n659_), .C1(new_n657_), .C2(new_n652_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  INV_X1    g462(.A(new_n310_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n626_), .A2(new_n306_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n310_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n306_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT47), .B(new_n665_), .C1(new_n666_), .C2(new_n306_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1330gat));
  NAND2_X1  g470(.A1(new_n389_), .A2(G50gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674_));
  AOI21_X1  g473(.A(G50gat), .B1(new_n626_), .B2(new_n389_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1331gat));
  NOR2_X1   g477(.A1(new_n484_), .A2(new_n524_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n543_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n597_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G57gat), .B1(new_n682_), .B2(new_n600_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n391_), .A2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n579_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n583_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n435_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n685_), .B2(new_n687_), .ZN(G1332gat));
  OAI21_X1  g487(.A(G64gat), .B1(new_n682_), .B2(new_n653_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT48), .ZN(new_n690_));
  INV_X1    g489(.A(new_n685_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n433_), .A3(new_n654_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1333gat));
  OR3_X1    g492(.A1(new_n685_), .A2(G71gat), .A3(new_n310_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n597_), .A2(new_n664_), .A3(new_n681_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(G71gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n682_), .B2(new_n269_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n691_), .A2(new_n442_), .A3(new_n389_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n684_), .A2(new_n625_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n402_), .B1(new_n705_), .B2(new_n583_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n643_), .A2(new_n644_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n680_), .A2(new_n542_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n330_), .A2(G85gat), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT112), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT113), .Z(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n709_), .B2(new_n653_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n705_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n403_), .A3(new_n604_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1337gat));
  AND3_X1   g516(.A1(new_n715_), .A2(new_n392_), .A3(new_n664_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n707_), .A2(new_n664_), .A3(new_n708_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G99gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n720_), .B(new_n722_), .ZN(G1338gat));
  NAND3_X1  g522(.A1(new_n715_), .A2(new_n393_), .A3(new_n389_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n389_), .B(new_n708_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n724_), .B(new_n730_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1339gat));
  NAND3_X1  g533(.A1(new_n504_), .A2(new_n510_), .A3(new_n507_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n505_), .B1(new_n512_), .B2(new_n506_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n520_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT116), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n735_), .A2(new_n739_), .A3(new_n520_), .A4(new_n736_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n523_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n478_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n466_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n454_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n467_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n468_), .A2(new_n422_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n469_), .B2(new_n426_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(KEYINPUT55), .A3(new_n456_), .A4(new_n454_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n746_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n475_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n475_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n742_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n572_), .B(new_n577_), .C1(new_n755_), .C2(KEYINPUT58), .ZN(new_n756_));
  INV_X1    g555(.A(new_n742_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n475_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n475_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n757_), .B(KEYINPUT58), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT117), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n755_), .B2(KEYINPUT58), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n756_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n524_), .A2(new_n478_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n479_), .A2(new_n741_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n575_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n524_), .A2(new_n478_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n767_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT57), .A3(new_n575_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n543_), .B1(new_n764_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n483_), .A2(new_n524_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n578_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n578_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  NOR4_X1   g584(.A1(new_n583_), .A2(new_n604_), .A3(new_n389_), .A4(new_n310_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n786_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT57), .B1(new_n774_), .B2(new_n575_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n770_), .B(new_n596_), .C1(new_n773_), .C2(new_n767_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n755_), .A2(KEYINPUT58), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n755_), .A2(new_n762_), .A3(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n760_), .A2(KEYINPUT117), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n642_), .A2(new_n794_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n542_), .B1(new_n793_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n578_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n780_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT118), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n777_), .A2(new_n802_), .A3(new_n783_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n790_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n787_), .B(new_n789_), .C1(new_n804_), .C2(new_n785_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n803_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n524_), .A3(new_n786_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n788_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n808_), .A3(KEYINPUT119), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1340gat));
  OAI21_X1  g612(.A(new_n787_), .B1(new_n804_), .B2(new_n785_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G120gat), .B1(new_n814_), .B2(new_n484_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n804_), .ZN(new_n816_));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n484_), .B2(KEYINPUT60), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(KEYINPUT60), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(KEYINPUT120), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT120), .B2(new_n818_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n816_), .B2(new_n821_), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n543_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n787_), .B(new_n824_), .C1(new_n804_), .C2(new_n785_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n806_), .A2(new_n542_), .A3(new_n786_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n804_), .A2(new_n833_), .A3(new_n596_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n642_), .B(new_n787_), .C1(new_n804_), .C2(new_n785_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n833_), .ZN(G1343gat));
  NAND3_X1  g636(.A1(new_n653_), .A2(new_n389_), .A3(new_n686_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n664_), .B(new_n838_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n524_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n483_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n839_), .B2(new_n542_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n838_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n806_), .A2(new_n310_), .A3(new_n542_), .A4(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n839_), .A2(new_n846_), .A3(new_n542_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n844_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1346gat));
  AOI21_X1  g654(.A(new_n664_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n596_), .A3(new_n848_), .ZN(new_n857_));
  INV_X1    g656(.A(G162gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n858_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n641_), .A2(new_n858_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n861_), .A2(new_n862_), .B1(new_n839_), .B2(new_n863_), .ZN(G1347gat));
  NAND3_X1  g663(.A1(new_n654_), .A2(new_n664_), .A3(new_n583_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT124), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n524_), .A3(new_n269_), .A4(new_n784_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT62), .B1(new_n867_), .B2(KEYINPUT22), .ZN(new_n868_));
  OAI21_X1  g667(.A(G169gat), .B1(new_n867_), .B2(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G169gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n868_), .ZN(G1348gat));
  AND3_X1   g671(.A1(new_n866_), .A2(new_n269_), .A3(new_n784_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G176gat), .B1(new_n873_), .B2(new_n483_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n806_), .A2(new_n269_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n806_), .A2(new_n877_), .A3(new_n269_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n876_), .A2(new_n866_), .A3(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n483_), .A2(G176gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n874_), .B1(new_n879_), .B2(new_n880_), .ZN(G1349gat));
  NAND4_X1  g680(.A1(new_n876_), .A2(new_n542_), .A3(new_n866_), .A4(new_n878_), .ZN(new_n882_));
  INV_X1    g681(.A(G183gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n543_), .A2(new_n283_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n882_), .A2(new_n883_), .B1(new_n873_), .B2(new_n884_), .ZN(G1350gat));
  NAND2_X1  g684(.A1(new_n873_), .A2(new_n642_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G190gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n873_), .A2(new_n341_), .A3(new_n596_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1351gat));
  NAND2_X1  g688(.A1(new_n654_), .A2(new_n373_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n856_), .A2(new_n524_), .A3(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g692(.A1(new_n856_), .A2(new_n483_), .A3(new_n891_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g694(.A(new_n543_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n856_), .A2(new_n891_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT126), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n897_), .B(new_n899_), .ZN(G1354gat));
  AND4_X1   g699(.A1(G218gat), .A2(new_n856_), .A3(new_n642_), .A4(new_n891_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n856_), .A2(new_n596_), .A3(new_n891_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n903_));
  AOI21_X1  g702(.A(G218gat), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n856_), .A2(new_n596_), .A3(new_n891_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT127), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n901_), .B1(new_n904_), .B2(new_n906_), .ZN(G1355gat));
endmodule


