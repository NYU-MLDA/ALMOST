//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n204_), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT87), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n210_), .A2(KEYINPUT21), .A3(new_n211_), .A4(new_n202_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT95), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT22), .B(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(KEYINPUT23), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(KEYINPUT24), .B2(new_n226_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n222_), .A2(KEYINPUT23), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT83), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n222_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n220_), .A2(new_n225_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n214_), .A2(new_n215_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n215_), .B1(new_n214_), .B2(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT20), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n220_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n228_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT25), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(new_n230_), .C1(new_n229_), .C2(new_n243_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n224_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n239_), .B1(new_n249_), .B2(new_n214_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n237_), .A2(new_n238_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT94), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT19), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n213_), .B(KEYINPUT90), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n236_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT20), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT97), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n249_), .A2(new_n214_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n257_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n255_), .B1(new_n264_), .B2(new_n254_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G64gat), .ZN(new_n268_));
  INV_X1    g067(.A(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n265_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G155gat), .B(G162gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT3), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT2), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n273_), .B1(new_n278_), .B2(KEYINPUT86), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(KEYINPUT86), .B2(new_n278_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n276_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n274_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n282_), .B(new_n283_), .C1(new_n273_), .C2(KEYINPUT1), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n284_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT84), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n292_), .A2(new_n303_), .A3(new_n296_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT96), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT96), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n305_), .B(new_n306_), .C1(new_n303_), .C2(new_n298_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n302_), .B1(new_n307_), .B2(new_n301_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT0), .ZN(new_n311_));
  INV_X1    g110(.A(G57gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(KEYINPUT98), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT98), .B1(new_n308_), .B2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n315_), .B2(new_n308_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n261_), .A2(new_n239_), .A3(new_n254_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n214_), .A2(new_n236_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n251_), .A2(new_n254_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n271_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n272_), .A2(new_n317_), .A3(new_n319_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n270_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n322_), .A2(new_n270_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n309_), .A2(KEYINPUT33), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n307_), .A2(new_n300_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n330_), .B(KEYINPUT33), .C1(new_n300_), .C2(new_n299_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n315_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n309_), .A2(KEYINPUT33), .A3(new_n316_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n248_), .B(KEYINPUT30), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT85), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n296_), .B(KEYINPUT31), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n342_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n341_), .B(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(new_n344_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n338_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n344_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n343_), .A2(new_n345_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n337_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G228gat), .ZN(new_n357_));
  INV_X1    g156(.A(G233gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n356_), .A2(new_n359_), .A3(new_n214_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n213_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(KEYINPUT89), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT89), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n355_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n360_), .B1(new_n366_), .B2(new_n359_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n367_), .A2(new_n371_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(new_n372_), .A2(new_n373_), .B1(new_n370_), .B2(new_n369_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n375_));
  XOR2_X1   g174(.A(G22gat), .B(G50gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT28), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n375_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n367_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n367_), .A2(new_n382_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .A4(new_n378_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT93), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n354_), .A2(new_n380_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n335_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n388_), .A3(new_n386_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n354_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n374_), .A2(new_n379_), .B1(new_n387_), .B2(KEYINPUT93), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n350_), .A2(new_n353_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n386_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT27), .B(new_n325_), .C1(new_n265_), .C2(new_n270_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n319_), .A2(new_n317_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n391_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT68), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G230gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT64), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G85gat), .A2(G92gat), .ZN(new_n407_));
  AND2_X1   g206(.A1(G85gat), .A2(G92gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(KEYINPUT9), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n269_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n314_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n409_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n416_), .A2(new_n417_), .A3(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n415_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n421_), .A3(new_n422_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT8), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n408_), .A2(new_n407_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n425_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G64gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G57gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n312_), .A2(G64gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT11), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT11), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G78gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(KEYINPUT11), .A3(new_n438_), .A4(new_n439_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n436_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n448_), .B(new_n425_), .C1(new_n435_), .C2(new_n434_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT12), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n436_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n406_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n406_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(KEYINPUT67), .A3(new_n406_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G120gat), .B(G148gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G204gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT5), .B(G176gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n404_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT67), .B1(new_n456_), .B2(new_n406_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n406_), .ZN(new_n468_));
  AOI211_X1 g267(.A(new_n458_), .B(new_n468_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n465_), .ZN(new_n471_));
  NOR4_X1   g270(.A1(new_n470_), .A2(KEYINPUT68), .A3(new_n455_), .A4(new_n471_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n466_), .A2(new_n472_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT13), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483_));
  INV_X1    g282(.A(G1gat), .ZN(new_n484_));
  INV_X1    g283(.A(G8gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT73), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G8gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n484_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n482_), .B(new_n483_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT73), .B(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n484_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n482_), .B1(new_n494_), .B2(new_n483_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n480_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n489_), .A2(new_n490_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n483_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n481_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n479_), .A3(new_n491_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G50gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G43gat), .ZN(new_n503_));
  INV_X1    g302(.A(G43gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G50gat), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n503_), .A2(new_n505_), .A3(KEYINPUT70), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT70), .B1(new_n503_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(G29gat), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(G50gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n502_), .A2(G43gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G29gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n503_), .A2(new_n505_), .A3(KEYINPUT70), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n508_), .A2(G36gat), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(G36gat), .B1(new_n508_), .B2(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G36gat), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n506_), .A2(new_n507_), .A3(G29gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n513_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n515_), .A3(G36gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n501_), .B1(new_n519_), .B2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n496_), .A2(new_n500_), .A3(new_n524_), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G169gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(G197gat), .Z(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT80), .ZN(new_n533_));
  INV_X1    g332(.A(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n523_), .A2(new_n524_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n501_), .A2(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n496_), .A2(new_n500_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n529_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n529_), .B2(new_n538_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n478_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n403_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n436_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n518_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n523_), .A2(KEYINPUT15), .A3(new_n524_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n436_), .B1(new_n519_), .B2(new_n525_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n535_), .A2(new_n436_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n556_), .A2(new_n560_), .A3(new_n554_), .A4(new_n549_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n562_), .A2(new_n567_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n571_), .B(new_n567_), .C1(new_n562_), .C2(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n549_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n556_), .B2(KEYINPUT71), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n553_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n568_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT72), .B1(new_n576_), .B2(new_n566_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n570_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT37), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n570_), .C1(new_n572_), .C2(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT78), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT78), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n501_), .A2(G231gat), .A3(G233gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n496_), .A2(new_n500_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n449_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n449_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n588_), .B(KEYINPUT17), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT79), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT79), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n600_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n583_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n544_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n399_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n484_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT38), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n578_), .B(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n402_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n389_), .B1(new_n324_), .B2(new_n334_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT101), .B(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n543_), .B(KEYINPUT99), .Z(new_n625_));
  NOR3_X1   g424(.A1(new_n624_), .A2(new_n609_), .A3(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n612_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n614_), .B1(new_n484_), .B2(new_n627_), .ZN(G1324gat));
  NAND2_X1  g427(.A1(new_n398_), .A2(new_n401_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n629_), .A3(new_n493_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n625_), .A2(new_n609_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n629_), .A3(new_n623_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n632_), .A2(new_n633_), .A3(G8gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n632_), .B2(G8gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n611_), .A2(new_n639_), .A3(new_n395_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n626_), .A2(new_n395_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n641_), .B2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(new_n392_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(G22gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT102), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n611_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n631_), .A2(new_n392_), .A3(new_n623_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G22gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n403_), .A2(KEYINPUT104), .A3(new_n656_), .A4(new_n583_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n583_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n656_), .B(new_n583_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n659_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n543_), .B(KEYINPUT99), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(new_n609_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(new_n665_), .A3(KEYINPUT44), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT44), .B1(new_n663_), .B2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n612_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT105), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n671_), .A3(new_n612_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(G29gat), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n616_), .A2(new_n608_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n544_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n513_), .A3(new_n612_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1328gat));
  NAND4_X1  g476(.A1(new_n544_), .A2(new_n520_), .A3(new_n629_), .A4(new_n674_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n629_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n666_), .A2(new_n667_), .A3(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(new_n520_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n685_));
  NOR2_X1   g484(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT107), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n685_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n663_), .A2(new_n665_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n663_), .A2(new_n665_), .A3(KEYINPUT44), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n629_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n680_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n685_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n688_), .A2(new_n697_), .ZN(G1329gat));
  AND3_X1   g497(.A1(new_n675_), .A2(new_n504_), .A3(new_n395_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n395_), .A3(new_n693_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G43gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n675_), .B2(new_n392_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n645_), .A2(new_n502_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n668_), .B2(new_n704_), .ZN(G1331gat));
  INV_X1    g504(.A(new_n478_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n541_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n403_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n610_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n312_), .A3(new_n612_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n608_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n624_), .A2(new_n399_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n712_), .B2(new_n312_), .ZN(G1332gat));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n437_), .A3(new_n629_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n624_), .A2(new_n711_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n437_), .B1(new_n715_), .B2(new_n629_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n709_), .A2(new_n721_), .A3(new_n395_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n624_), .A2(new_n354_), .A3(new_n711_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n723_), .A2(KEYINPUT108), .A3(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT108), .B1(new_n723_), .B2(new_n721_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(KEYINPUT49), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT49), .B1(new_n724_), .B2(new_n725_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n726_), .B2(new_n727_), .ZN(G1334gat));
  INV_X1    g527(.A(G78gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n709_), .A2(new_n729_), .A3(new_n392_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n645_), .B(new_n711_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(new_n731_), .B2(new_n729_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n623_), .A2(new_n392_), .A3(new_n608_), .A4(new_n707_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(G78gat), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n732_), .A2(new_n735_), .A3(KEYINPUT50), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT50), .B1(new_n732_), .B2(new_n735_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n730_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT110), .B(new_n730_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NAND3_X1  g541(.A1(new_n663_), .A2(new_n609_), .A3(new_n707_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n399_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n708_), .A2(new_n674_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n314_), .A3(new_n612_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1336gat));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n629_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n269_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n411_), .A2(new_n412_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n629_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n745_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT112), .B(new_n751_), .C1(new_n745_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n743_), .B2(new_n354_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n354_), .A2(new_n417_), .A3(new_n416_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n747_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n428_), .B1(new_n764_), .B2(KEYINPUT52), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n743_), .B2(new_n645_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(KEYINPUT113), .A3(new_n767_), .ZN(new_n768_));
  OAI221_X1 g567(.A(new_n765_), .B1(new_n764_), .B2(KEYINPUT52), .C1(new_n743_), .C2(new_n645_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n747_), .A2(new_n428_), .A3(new_n392_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n768_), .A2(new_n773_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  OAI21_X1  g574(.A(new_n541_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT115), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n452_), .A2(new_n454_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n468_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n465_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT68), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n461_), .A2(new_n404_), .A3(new_n465_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n541_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n455_), .B(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n452_), .A2(new_n406_), .A3(new_n454_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n452_), .A2(KEYINPUT116), .A3(new_n406_), .A4(new_n454_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n465_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n786_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n779_), .A2(new_n787_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n455_), .A2(KEYINPUT55), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n471_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n777_), .A2(new_n785_), .A3(new_n796_), .A4(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n526_), .A2(new_n527_), .A3(new_n534_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n528_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(new_n532_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n529_), .A2(new_n538_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n532_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n473_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n802_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n616_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n800_), .A2(new_n786_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n471_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n806_), .A2(new_n808_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n582_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n819_), .A3(new_n815_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n812_), .A2(new_n813_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n811_), .A2(new_n616_), .A3(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n608_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n608_), .B2(new_n542_), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT114), .B(new_n541_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n474_), .A4(new_n582_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n474_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n832_), .B2(new_n583_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n810_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n783_), .A2(new_n784_), .A3(new_n541_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n784_), .B1(new_n783_), .B2(new_n541_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n796_), .A2(new_n801_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n836_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n578_), .B(KEYINPUT100), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n813_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n821_), .A2(new_n822_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n824_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n609_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n831_), .A2(new_n833_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n396_), .A2(new_n629_), .A3(new_n399_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n835_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n541_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  INV_X1    g655(.A(new_n824_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n823_), .B2(KEYINPUT120), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n843_), .A2(new_n844_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n608_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n856_), .B(new_n850_), .C1(new_n862_), .C2(new_n834_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT121), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n855_), .A2(new_n866_), .A3(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n542_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n854_), .B1(new_n868_), .B2(new_n853_), .ZN(G1340gat));
  NOR2_X1   g668(.A1(new_n706_), .A2(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n852_), .B1(KEYINPUT60), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n478_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G120gat), .B1(new_n872_), .B2(new_n864_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n852_), .A2(new_n875_), .A3(new_n608_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n609_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1342gat));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n852_), .A2(new_n879_), .A3(new_n842_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n582_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT122), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n884_), .B(new_n880_), .C1(new_n881_), .C2(new_n879_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1343gat));
  AND2_X1   g685(.A1(new_n835_), .A2(new_n849_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n395_), .B1(new_n394_), .B2(new_n386_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n887_), .A2(new_n612_), .A3(new_n888_), .A4(new_n682_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n542_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n706_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n609_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n889_), .B2(new_n582_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n616_), .A2(G162gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n889_), .B2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n682_), .A2(new_n612_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n395_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n542_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT123), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n645_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n862_), .A2(new_n834_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G169gat), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT62), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n392_), .A3(new_n901_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n218_), .A3(new_n541_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n908_), .B2(new_n478_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n887_), .A2(new_n645_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n901_), .A2(new_n219_), .A3(new_n706_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  INV_X1    g713(.A(new_n908_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n915_), .A2(new_n229_), .A3(new_n609_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n912_), .A2(new_n395_), .A3(new_n608_), .A4(new_n900_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n917_), .B2(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n916_), .B1(new_n919_), .B2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n915_), .B2(new_n582_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n908_), .A2(new_n842_), .A3(new_n230_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  NAND4_X1  g723(.A1(new_n835_), .A2(new_n849_), .A3(new_n888_), .A4(new_n900_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT125), .Z(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n541_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT126), .B(G197gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n478_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g730(.A(new_n609_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n926_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  XOR2_X1   g733(.A(new_n933_), .B(new_n934_), .Z(G1354gat));
  NOR2_X1   g734(.A1(new_n616_), .A2(G218gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n926_), .A2(new_n936_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n926_), .A2(new_n583_), .ZN(new_n938_));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  OAI211_X1 g738(.A(KEYINPUT127), .B(new_n937_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  INV_X1    g740(.A(new_n937_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n939_), .B1(new_n926_), .B2(new_n583_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n944_), .ZN(G1355gat));
endmodule


