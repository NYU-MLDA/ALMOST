//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT88), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT90), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT89), .B1(new_n217_), .B2(KEYINPUT22), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n218_), .C1(new_n219_), .C2(KEYINPUT89), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n212_), .A3(new_n215_), .A4(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n204_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n205_), .A2(KEYINPUT86), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n225_), .B(KEYINPUT25), .Z(new_n226_));
  NOR3_X1   g025(.A1(new_n206_), .A2(KEYINPUT87), .A3(KEYINPUT26), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(KEYINPUT87), .ZN(new_n229_));
  OAI221_X1 g028(.A(new_n223_), .B1(new_n224_), .B2(new_n211_), .C1(new_n226_), .C2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT30), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G15gat), .B(G43gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n232_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n233_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n232_), .A2(KEYINPUT92), .A3(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G127gat), .B(G134gat), .ZN(new_n248_));
  INV_X1    g047(.A(G120gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT93), .B(G113gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT31), .ZN(new_n253_));
  OR4_X1    g052(.A1(KEYINPUT94), .A2(new_n242_), .A3(new_n247_), .A4(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT94), .B1(new_n242_), .B2(new_n247_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n241_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n258_), .A3(new_n253_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT95), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT98), .ZN(new_n265_));
  INV_X1    g064(.A(G141gat), .ZN(new_n266_));
  INV_X1    g065(.A(G148gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OR3_X1    g067(.A1(new_n268_), .A2(KEYINPUT96), .A3(KEYINPUT3), .ZN(new_n269_));
  NAND2_X1  g068(.A1(KEYINPUT97), .A2(KEYINPUT2), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(KEYINPUT97), .A2(KEYINPUT2), .ZN(new_n272_));
  OAI211_X1 g071(.A(G141gat), .B(G148gat), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n274_), .A2(new_n270_), .B1(KEYINPUT96), .B2(KEYINPUT3), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n268_), .B1(KEYINPUT96), .B2(KEYINPUT3), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n269_), .A2(new_n273_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT98), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n262_), .A2(new_n278_), .A3(new_n263_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n265_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n262_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n263_), .B(KEYINPUT1), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n268_), .B(new_n274_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT100), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G228gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT101), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(new_n291_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT100), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n287_), .A2(new_n289_), .A3(new_n298_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n289_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n298_), .B(KEYINPUT102), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(new_n300_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT103), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n302_), .A2(new_n305_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n306_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT103), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n280_), .A2(new_n299_), .A3(new_n283_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G22gat), .B(G50gat), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT99), .B(KEYINPUT28), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n317_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n318_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n310_), .A2(new_n315_), .A3(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n313_), .A2(new_n324_), .A3(new_n314_), .A4(new_n307_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n296_), .A2(new_n297_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT102), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT102), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n298_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n207_), .A2(new_n211_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n219_), .A2(new_n216_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT104), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n228_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n224_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n210_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n223_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n330_), .A2(new_n332_), .A3(new_n335_), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n231_), .B2(new_n298_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT19), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n329_), .A2(new_n221_), .A3(new_n230_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(KEYINPUT105), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT105), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n339_), .A2(new_n352_), .A3(new_n223_), .A4(new_n341_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n351_), .A2(new_n353_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT20), .B(new_n350_), .C1(new_n354_), .C2(new_n329_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n349_), .B1(new_n355_), .B2(new_n348_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT18), .B(G64gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n348_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n354_), .A2(new_n329_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n348_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n345_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n366_), .A3(new_n360_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n362_), .A2(KEYINPUT27), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n366_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n361_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT27), .B1(new_n370_), .B2(new_n367_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT110), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  INV_X1    g173(.A(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n284_), .A2(KEYINPUT106), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT106), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n280_), .A2(new_n383_), .A3(new_n283_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n384_), .A3(new_n252_), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n250_), .B(new_n251_), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n284_), .A2(KEYINPUT106), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n284_), .A2(new_n381_), .A3(new_n252_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n380_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n378_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n391_), .A3(new_n378_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n328_), .A2(new_n372_), .A3(new_n373_), .A4(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n326_), .A2(new_n394_), .A3(new_n393_), .A4(new_n327_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n362_), .A2(KEYINPUT27), .A3(new_n367_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n367_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n360_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n399_), .B1(new_n402_), .B2(KEYINPUT27), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT110), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n370_), .A2(new_n367_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n388_), .A2(new_n380_), .A3(new_n389_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT108), .ZN(new_n408_));
  INV_X1    g207(.A(new_n378_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n385_), .A2(new_n387_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT107), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n411_), .B2(new_n380_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n406_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n392_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n363_), .A2(new_n366_), .A3(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT109), .Z(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n393_), .A2(new_n394_), .B1(new_n356_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n328_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n260_), .B1(new_n405_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n254_), .A2(new_n396_), .A3(new_n259_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n328_), .A2(new_n403_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G57gat), .B(G64gat), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT67), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G71gat), .ZN(new_n434_));
  INV_X1    g233(.A(G78gat), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT11), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n433_), .A2(G71gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n431_), .A2(KEYINPUT67), .ZN(new_n441_));
  OAI21_X1  g240(.A(G78gat), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT11), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n430_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(KEYINPUT11), .A3(new_n443_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n430_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n438_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n451_), .B2(new_n447_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n436_), .A2(new_n437_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n430_), .B1(new_n453_), .B2(KEYINPUT11), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT68), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G92gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT64), .B1(new_n375_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT9), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT64), .B(new_n460_), .C1(new_n375_), .C2(new_n457_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n459_), .B(new_n461_), .C1(G85gat), .C2(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(KEYINPUT10), .B(G99gat), .Z(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(KEYINPUT66), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n464_), .A2(new_n466_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G85gat), .B(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n472_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n467_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n472_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n471_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n456_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n452_), .A2(new_n454_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n498_), .A2(new_n494_), .A3(new_n491_), .A4(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G120gat), .B(G148gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT72), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G176gat), .B(G204gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT70), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n496_), .A2(new_n502_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT13), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT79), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G1gat), .B(G8gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G29gat), .ZN(new_n526_));
  INV_X1    g325(.A(G36gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G50gat), .ZN(new_n531_));
  INV_X1    g330(.A(G50gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n532_), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT73), .B(G43gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n535_), .A3(new_n533_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n525_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT15), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n531_), .A2(new_n535_), .A3(new_n533_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n535_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n537_), .A2(KEYINPUT15), .A3(new_n538_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n525_), .A2(KEYINPUT84), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n525_), .A2(new_n539_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT84), .B1(new_n525_), .B2(new_n549_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n550_), .A2(new_n542_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G169gat), .B(G197gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT85), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n554_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n515_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n547_), .A2(new_n548_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n489_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT75), .B1(new_n565_), .B2(KEYINPUT35), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n539_), .B(new_n471_), .C1(new_n483_), .C2(new_n488_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n565_), .A2(KEYINPUT75), .A3(KEYINPUT35), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n563_), .A2(new_n566_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n567_), .A2(KEYINPUT74), .A3(new_n566_), .A4(new_n568_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(KEYINPUT35), .A3(new_n565_), .A4(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(KEYINPUT35), .A3(new_n565_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n567_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n563_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT76), .B(G190gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT36), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n571_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n583_), .B2(KEYINPUT77), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n525_), .B(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(new_n500_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT17), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT81), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n500_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n594_), .A2(new_n456_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n594_), .A2(new_n456_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n600_), .A2(KEYINPUT17), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT82), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n592_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT83), .Z(new_n613_));
  AND3_X1   g412(.A1(new_n429_), .A2(new_n561_), .A3(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n519_), .A3(new_n395_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT38), .ZN(new_n616_));
  INV_X1    g415(.A(new_n611_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT113), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n413_), .A2(new_n415_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n397_), .B(new_n404_), .C1(new_n619_), .C2(new_n328_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n620_), .A2(new_n260_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT112), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n571_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n580_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n622_), .B(new_n585_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n618_), .B1(new_n621_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n429_), .A2(KEYINPUT113), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n617_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n561_), .B(KEYINPUT111), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n395_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G1gat), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n616_), .A2(new_n635_), .ZN(G1324gat));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n631_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n637_), .A2(new_n633_), .A3(new_n611_), .A4(new_n403_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT114), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT114), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(G8gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(KEYINPUT39), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n614_), .A2(new_n520_), .A3(new_n403_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n639_), .A2(KEYINPUT114), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n643_), .A2(KEYINPUT40), .A3(new_n644_), .A4(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n260_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n614_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n632_), .A2(new_n633_), .A3(new_n653_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n655_), .B2(G15gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n614_), .A2(new_n659_), .A3(new_n328_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n632_), .A2(new_n633_), .A3(new_n328_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G22gat), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1327gat));
  NAND3_X1  g464(.A1(new_n429_), .A2(new_n617_), .A3(new_n628_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n666_), .A2(new_n560_), .A3(new_n515_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n395_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n621_), .B2(new_n592_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n592_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n429_), .A2(KEYINPUT43), .A3(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n670_), .A2(new_n672_), .A3(new_n633_), .A4(new_n617_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n526_), .B(new_n396_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n668_), .B1(new_n675_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n667_), .A2(new_n527_), .A3(new_n403_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n372_), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n673_), .A2(new_n674_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n527_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n679_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n681_), .A3(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1329gat));
  NAND4_X1  g488(.A1(new_n677_), .A2(G43gat), .A3(new_n653_), .A4(new_n684_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n667_), .A2(new_n653_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(G43gat), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n667_), .B2(new_n328_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n677_), .A2(G50gat), .A3(new_n684_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n328_), .ZN(G1331gat));
  INV_X1    g495(.A(new_n515_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n559_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n632_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT116), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT116), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n632_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n702_));
  AND4_X1   g501(.A1(G57gat), .A2(new_n700_), .A3(new_n395_), .A4(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n613_), .A2(new_n515_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(KEYINPUT115), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n559_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n621_), .B1(new_n704_), .B2(KEYINPUT115), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n395_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n703_), .A2(new_n710_), .ZN(G1332gat));
  OR3_X1    g510(.A1(new_n708_), .A2(G64gat), .A3(new_n372_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(new_n403_), .A3(new_n702_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1333gat));
  NAND3_X1  g516(.A1(new_n709_), .A2(new_n431_), .A3(new_n653_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n700_), .A2(new_n653_), .A3(new_n702_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G71gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G71gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  NAND3_X1  g522(.A1(new_n709_), .A2(new_n435_), .A3(new_n328_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n700_), .A2(new_n328_), .A3(new_n702_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1335gat));
  AND2_X1   g528(.A1(new_n670_), .A2(new_n672_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n617_), .A3(new_n698_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n396_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n666_), .A2(new_n559_), .A3(new_n697_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n375_), .A3(new_n395_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT117), .Z(G1336gat));
  NOR3_X1   g535(.A1(new_n731_), .A2(new_n457_), .A3(new_n372_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G92gat), .B1(new_n733_), .B2(new_n403_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1337gat));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n468_), .A3(new_n653_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT118), .ZN(new_n741_));
  INV_X1    g540(.A(G99gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n731_), .A2(new_n260_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n741_), .B(new_n745_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n733_), .A2(new_n469_), .A3(new_n328_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n730_), .A2(new_n617_), .A3(new_n328_), .A4(new_n698_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(G106gat), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n751_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n750_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n427_), .A2(new_n395_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n502_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n480_), .A2(new_n482_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT8), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n499_), .B1(new_n769_), .B2(new_n471_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n770_), .A2(KEYINPUT12), .B1(new_n456_), .B2(new_n490_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(KEYINPUT55), .A3(new_n494_), .A4(new_n498_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n765_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n498_), .A2(new_n491_), .A3(new_n501_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n495_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(new_n495_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n773_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n508_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(G229gat), .A3(G233gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n541_), .A2(new_n542_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n557_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n554_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n557_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n496_), .A2(new_n502_), .A3(new_n779_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  INV_X1    g587(.A(new_n777_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n774_), .A2(new_n775_), .A3(new_n495_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n788_), .B(new_n508_), .C1(new_n791_), .C2(new_n773_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n780_), .A2(new_n786_), .A3(new_n787_), .A4(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n780_), .A2(new_n559_), .A3(new_n787_), .A4(new_n792_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n786_), .B1(new_n511_), .B2(new_n510_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n630_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n798_), .A2(new_n671_), .B1(new_n799_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n628_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT122), .B1(new_n805_), .B2(KEYINPUT57), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n611_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n697_), .A2(new_n592_), .A3(new_n611_), .A4(new_n560_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n653_), .B(new_n763_), .C1(new_n809_), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n793_), .A2(new_n794_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n671_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n799_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n805_), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(new_n824_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n812_), .B1(new_n827_), .B2(new_n617_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(new_n260_), .A3(new_n762_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n814_), .B1(new_n828_), .B2(KEYINPUT123), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n817_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n761_), .B1(new_n832_), .B2(new_n559_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n559_), .A2(new_n761_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n813_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT124), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n560_), .B1(new_n817_), .B2(new_n831_), .ZN(new_n838_));
  OAI221_X1 g637(.A(new_n837_), .B1(new_n813_), .B2(new_n834_), .C1(new_n838_), .C2(new_n761_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1340gat));
  NOR2_X1   g639(.A1(new_n697_), .A2(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n829_), .B1(KEYINPUT60), .B2(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n832_), .A2(new_n515_), .A3(new_n842_), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n843_), .A2(new_n249_), .B1(KEYINPUT60), .B2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n829_), .B2(new_n611_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n832_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n617_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n829_), .B2(new_n628_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n846_), .A2(new_n592_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g650(.A(new_n828_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n260_), .A2(new_n395_), .A3(new_n328_), .A4(new_n372_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT125), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n560_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n266_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n697_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n267_), .ZN(G1345gat));
  NOR2_X1   g658(.A1(new_n855_), .A2(new_n617_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT61), .B(G155gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  INV_X1    g661(.A(G162gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n855_), .A2(new_n863_), .A3(new_n592_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n852_), .A2(new_n628_), .A3(new_n854_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n328_), .A2(new_n372_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n852_), .A2(new_n426_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n560_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n867_), .B1(new_n870_), .B2(new_n217_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n219_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT62), .B(G169gat), .C1(new_n869_), .C2(new_n560_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(G1348gat));
  NOR2_X1   g673(.A1(new_n869_), .A2(new_n697_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n216_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n869_), .A2(new_n617_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n338_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n205_), .B2(new_n877_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n869_), .B2(new_n592_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n628_), .A2(new_n228_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n869_), .B2(new_n881_), .ZN(G1351gat));
  INV_X1    g681(.A(new_n398_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n653_), .A2(new_n372_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n852_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n559_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n515_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g689(.A1(new_n885_), .A2(new_n617_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n892_));
  INV_X1    g691(.A(G211gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n891_), .A2(new_n898_), .A3(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n892_), .A2(new_n893_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n897_), .A2(new_n892_), .A3(new_n899_), .A4(new_n893_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1354gat));
  NAND3_X1  g703(.A1(new_n886_), .A2(G218gat), .A3(new_n671_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n885_), .A2(new_n630_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(G218gat), .B2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


