//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT82), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT82), .A4(new_n207_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n215_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n217_), .B1(new_n220_), .B2(KEYINPUT23), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT80), .B(G183gat), .Z(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n216_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(KEYINPUT23), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n218_), .B(KEYINPUT81), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(KEYINPUT23), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(G169gat), .B(G176gat), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT24), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n222_), .B2(KEYINPUT25), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT26), .B(G190gat), .Z(new_n235_));
  OAI211_X1 g034(.A(new_n229_), .B(new_n232_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n225_), .A2(new_n226_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n226_), .B1(new_n225_), .B2(new_n236_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  INV_X1    g039(.A(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G127gat), .B(G134gat), .Z(new_n244_));
  XOR2_X1   g043(.A(G113gat), .B(G120gat), .Z(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT85), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  XOR2_X1   g047(.A(new_n243_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n243_), .B(new_n248_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G211gat), .B(G218gat), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT91), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(G204gat), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n266_), .C1(G197gat), .C2(new_n265_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n261_), .A2(KEYINPUT21), .A3(new_n267_), .A4(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT92), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n260_), .B2(KEYINPUT91), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n275_), .A2(KEYINPUT92), .A3(new_n267_), .A4(new_n270_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n263_), .A2(G204gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n265_), .A2(G197gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT21), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n268_), .C1(new_n267_), .C2(KEYINPUT21), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT88), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT86), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT3), .ZN(new_n292_));
  OR3_X1    g091(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n292_), .B(new_n293_), .C1(new_n289_), .C2(new_n287_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n285_), .B(new_n286_), .C1(new_n290_), .C2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n291_), .B(KEYINPUT87), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n286_), .B(KEYINPUT1), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n296_), .B(new_n288_), .C1(new_n284_), .C2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n282_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G78gat), .B(G106gat), .Z(new_n302_));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n305_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n300_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT28), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n311_), .A2(new_n307_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G22gat), .B(G50gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n295_), .A2(new_n298_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT4), .B1(new_n248_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n248_), .A2(new_n322_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n244_), .A2(new_n245_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n295_), .B(new_n298_), .C1(new_n247_), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n327_), .B2(KEYINPUT4), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT98), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n332_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT19), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n225_), .A2(new_n236_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT84), .ZN(new_n348_));
  INV_X1    g147(.A(new_n282_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n225_), .A2(new_n226_), .A3(new_n236_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n354_));
  MUX2_X1   g153(.A(new_n231_), .B(new_n353_), .S(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n235_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT25), .B(G183gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n229_), .B1(G183gat), .B2(G190gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n211_), .B(KEYINPUT95), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n204_), .A2(new_n206_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n207_), .B2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n358_), .A2(new_n221_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n349_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n352_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT93), .B1(new_n351_), .B2(KEYINPUT20), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n346_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n349_), .B2(new_n363_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n282_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n346_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT97), .ZN(new_n376_));
  XOR2_X1   g175(.A(G64gat), .B(G92gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n344_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT93), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n237_), .A2(new_n238_), .A3(new_n282_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n368_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n346_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n364_), .A4(new_n352_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n346_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n390_), .A2(KEYINPUT99), .A3(new_n382_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT99), .B1(new_n390_), .B2(new_n382_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n383_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n367_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n380_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n374_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n328_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n329_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n339_), .B1(new_n333_), .B2(new_n330_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT33), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n342_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n341_), .A2(KEYINPUT33), .ZN(new_n403_));
  AND4_X1   g202(.A1(new_n394_), .A2(new_n396_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n321_), .B1(new_n393_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n321_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n390_), .A2(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT100), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT100), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n390_), .A2(new_n409_), .A3(new_n395_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n386_), .A2(new_n364_), .A3(new_n352_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n372_), .B1(new_n412_), .B2(new_n346_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n413_), .B2(new_n380_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n344_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n394_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n380_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n406_), .A2(new_n415_), .A3(new_n416_), .A4(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n259_), .B1(new_n405_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n319_), .A2(new_n344_), .A3(new_n320_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n259_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n415_), .A2(KEYINPUT101), .A3(new_n419_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT101), .B1(new_n415_), .B2(new_n419_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT102), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n394_), .A2(KEYINPUT27), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n409_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n432_));
  AOI211_X1 g231(.A(KEYINPUT100), .B(new_n380_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT27), .B1(new_n396_), .B2(new_n394_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n430_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n415_), .A2(new_n419_), .A3(KEYINPUT101), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(KEYINPUT102), .A3(new_n424_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n421_), .B1(new_n429_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G190gat), .B(G218gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT73), .ZN(new_n442_));
  XOR2_X1   g241(.A(G134gat), .B(G162gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT36), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G106gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  OAI22_X1  g251(.A1(new_n452_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  OR4_X1    g252(.A1(new_n452_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n449_), .A2(new_n451_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT8), .B1(new_n458_), .B2(KEYINPUT67), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT64), .B(G106gat), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT10), .B(G99gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n465_), .A2(new_n449_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n456_), .A2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n451_), .A2(new_n469_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n459_), .A2(new_n460_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n459_), .A2(new_n460_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G29gat), .B(G36gat), .Z(new_n474_));
  XOR2_X1   g273(.A(G43gat), .B(G50gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G232gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT34), .ZN(new_n479_));
  OAI22_X1  g278(.A1(new_n473_), .A2(new_n477_), .B1(KEYINPUT35), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n476_), .B(KEYINPUT15), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n473_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(KEYINPUT35), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n484_), .A2(KEYINPUT36), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n445_), .B1(new_n485_), .B2(new_n444_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n484_), .A2(KEYINPUT74), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT68), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(KEYINPUT11), .B2(new_n492_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  INV_X1    g301(.A(G8gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n501_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513_));
  XOR2_X1   g312(.A(G127gat), .B(G155gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT16), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n512_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n501_), .B2(new_n511_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n499_), .B(KEYINPUT75), .ZN(new_n520_));
  INV_X1    g319(.A(new_n511_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n517_), .B(KEYINPUT17), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n440_), .A2(new_n491_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n499_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT12), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n473_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT12), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n501_), .A2(KEYINPUT70), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT70), .B1(new_n501_), .B2(new_n534_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n531_), .B(new_n532_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n530_), .B2(new_n528_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G120gat), .B(G148gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G176gat), .B(G204gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT71), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n540_), .B(new_n546_), .Z(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT13), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n476_), .A2(new_n508_), .A3(new_n507_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT76), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n477_), .A2(new_n509_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT77), .Z(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n481_), .A2(new_n509_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n555_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT78), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n557_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n560_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n563_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n567_), .A2(KEYINPUT79), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(KEYINPUT79), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n549_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n527_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n202_), .B1(new_n573_), .B2(new_n344_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT103), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n440_), .A2(new_n571_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n526_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n488_), .A2(KEYINPUT37), .A3(new_n489_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT37), .B1(new_n488_), .B2(new_n489_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND4_X1   g379(.A1(new_n548_), .A2(new_n576_), .A3(new_n577_), .A4(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n202_), .A3(new_n344_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT38), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n575_), .A2(new_n583_), .ZN(G1324gat));
  INV_X1    g383(.A(new_n438_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n503_), .B1(new_n573_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT39), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n503_), .A3(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT40), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(G1325gat));
  AOI21_X1  g390(.A(new_n251_), .B1(new_n573_), .B2(new_n259_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT41), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n581_), .A2(new_n251_), .A3(new_n259_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(G1326gat));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n573_), .B2(new_n406_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT42), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n581_), .A2(new_n596_), .A3(new_n406_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1327gat));
  NAND2_X1  g399(.A1(new_n491_), .A2(new_n526_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n549_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n576_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(G29gat), .B1(new_n603_), .B2(new_n344_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT43), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n440_), .B2(new_n580_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n405_), .A2(new_n420_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n259_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT102), .B1(new_n438_), .B2(new_n424_), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n428_), .B(new_n423_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n579_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n488_), .A2(KEYINPUT37), .A3(new_n489_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(KEYINPUT43), .A3(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n606_), .A2(new_n616_), .A3(new_n572_), .A4(new_n526_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  AND4_X1   g422(.A1(new_n572_), .A2(new_n606_), .A3(new_n526_), .A4(new_n616_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT44), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n344_), .A2(G29gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n604_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n617_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n621_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n585_), .B(new_n625_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  INV_X1    g433(.A(G36gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n438_), .B(KEYINPUT105), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n603_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n630_), .B1(new_n634_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1329gat));
  INV_X1    g441(.A(new_n603_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n241_), .B1(new_n643_), .B2(new_n608_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n259_), .A2(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n626_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1330gat));
  INV_X1    g447(.A(G50gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n406_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT109), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n603_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n406_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n649_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n321_), .B1(new_n624_), .B2(KEYINPUT44), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n632_), .B2(new_n631_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT108), .B1(new_n658_), .B2(G50gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n652_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT110), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT110), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n662_), .B(new_n652_), .C1(new_n656_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1331gat));
  NOR3_X1   g463(.A1(new_n615_), .A2(new_n548_), .A3(new_n526_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n440_), .A2(new_n570_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n344_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n548_), .A2(new_n570_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n527_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n344_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(new_n669_), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n672_), .B2(new_n637_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NOR2_X1   g476(.A1(new_n636_), .A2(G64gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT111), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n667_), .B2(new_n679_), .ZN(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n672_), .B2(new_n259_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT49), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n259_), .A2(new_n681_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT112), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n668_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT113), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n672_), .B2(new_n406_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT50), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n668_), .A2(new_n690_), .A3(new_n406_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1335gat));
  NOR4_X1   g493(.A1(new_n440_), .A2(new_n601_), .A3(new_n570_), .A4(new_n548_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G85gat), .B1(new_n695_), .B2(new_n344_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n606_), .A2(new_n526_), .A3(new_n616_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n671_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n344_), .A2(G85gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT114), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n699_), .B2(new_n701_), .ZN(G1336gat));
  OAI21_X1  g501(.A(G92gat), .B1(new_n698_), .B2(new_n636_), .ZN(new_n703_));
  INV_X1    g502(.A(G92gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n695_), .A2(new_n704_), .A3(new_n585_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1337gat));
  OAI21_X1  g505(.A(G99gat), .B1(new_n698_), .B2(new_n608_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n695_), .A2(new_n464_), .A3(new_n259_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g509(.A1(new_n695_), .A2(new_n462_), .A3(new_n406_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n699_), .A2(new_n406_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n448_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT53), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT53), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n711_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1339gat));
  NAND4_X1  g521(.A1(new_n580_), .A2(new_n571_), .A3(new_n548_), .A4(new_n577_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT54), .Z(new_n724_));
  OR2_X1    g523(.A1(new_n568_), .A2(new_n569_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n559_), .A2(new_n555_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n563_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n537_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n531_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n538_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(KEYINPUT55), .A3(new_n537_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n732_), .A2(KEYINPUT55), .A3(new_n538_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT116), .ZN(new_n737_));
  INV_X1    g536(.A(new_n545_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n735_), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(KEYINPUT119), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT119), .B1(new_n741_), .B2(new_n742_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n738_), .A4(new_n740_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT118), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n731_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT120), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT58), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT119), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n734_), .A2(new_n735_), .A3(new_n739_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n739_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n545_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n754_), .B2(KEYINPUT56), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n746_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n741_), .A2(KEYINPUT119), .A3(new_n742_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n755_), .A2(new_n756_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n731_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(KEYINPUT120), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n750_), .A2(new_n615_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n570_), .A2(new_n730_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n753_), .A2(new_n545_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n740_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n746_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n725_), .A2(new_n728_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(new_n547_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n491_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(KEYINPUT57), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n741_), .A2(new_n742_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n766_), .B1(new_n778_), .B2(new_n746_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n772_), .A2(new_n547_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n490_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n777_), .B1(new_n781_), .B2(KEYINPUT117), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n776_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n765_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n724_), .B1(new_n784_), .B2(new_n526_), .ZN(new_n785_));
  NOR4_X1   g584(.A1(new_n585_), .A2(new_n416_), .A3(new_n608_), .A4(new_n406_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n570_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT59), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n577_), .B1(new_n765_), .B2(new_n783_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT59), .B(new_n786_), .C1(new_n792_), .C2(new_n724_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n570_), .A2(G113gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT121), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n789_), .B1(new_n794_), .B2(new_n796_), .ZN(G1340gat));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n788_), .B(new_n799_), .C1(KEYINPUT60), .C2(new_n798_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n548_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n798_), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(new_n803_), .A3(new_n577_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n526_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1342gat));
  XNOR2_X1  g605(.A(KEYINPUT122), .B(G134gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n615_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n724_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n774_), .B2(new_n775_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n781_), .A2(KEYINPUT117), .A3(new_n777_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n762_), .A2(KEYINPUT120), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n580_), .B1(new_n814_), .B2(KEYINPUT58), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n764_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n810_), .B1(new_n816_), .B2(new_n577_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT59), .B1(new_n817_), .B2(new_n786_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n793_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n809_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n491_), .B(new_n786_), .C1(new_n792_), .C2(new_n724_), .ZN(new_n822_));
  INV_X1    g621(.A(G134gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n821_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n808_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n824_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT123), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1343gat));
  NOR2_X1   g628(.A1(new_n259_), .A2(new_n321_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n636_), .A2(new_n344_), .A3(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n785_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n570_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n549_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n577_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  INV_X1    g638(.A(G162gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n840_), .A3(new_n491_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(new_n615_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n840_), .ZN(G1347gat));
  OAI211_X1 g643(.A(new_n424_), .B(new_n637_), .C1(new_n792_), .C2(new_n724_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G169gat), .B1(new_n845_), .B2(new_n571_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n845_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n570_), .A3(new_n361_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n849_), .A3(new_n851_), .ZN(G1348gat));
  NOR2_X1   g651(.A1(new_n845_), .A2(new_n548_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n207_), .ZN(G1349gat));
  NOR2_X1   g653(.A1(new_n845_), .A2(new_n526_), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n222_), .B(new_n357_), .S(new_n855_), .Z(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n845_), .B2(new_n580_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n490_), .A2(new_n235_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n845_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n857_), .B(KEYINPUT124), .C1(new_n845_), .C2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1351gat));
  NAND2_X1  g663(.A1(new_n830_), .A2(new_n416_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT125), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n637_), .B(new_n866_), .C1(new_n792_), .C2(new_n724_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n571_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n263_), .A2(KEYINPUT126), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n263_), .A2(KEYINPUT126), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n868_), .B2(new_n870_), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n867_), .A2(new_n548_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n265_), .ZN(G1353gat));
  NOR2_X1   g673(.A1(new_n867_), .A2(new_n526_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT63), .B(G211gat), .Z(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(G1354gat));
  OAI21_X1  g677(.A(G218gat), .B1(new_n867_), .B2(new_n580_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n490_), .A2(G218gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n867_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT127), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n879_), .B(new_n884_), .C1(new_n867_), .C2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1355gat));
endmodule


