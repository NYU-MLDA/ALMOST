//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT19), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G218gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G211gat), .ZN(new_n210_));
  INV_X1    g009(.A(G211gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G218gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n215_));
  AND2_X1   g014(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(G204gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(G197gat), .B2(G204gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n214_), .A2(new_n215_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(G204gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G197gat), .A2(G204gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT21), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n210_), .A2(new_n212_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT92), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n223_), .A2(KEYINPUT21), .A3(new_n225_), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n222_), .A2(new_n226_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT101), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n234_), .A2(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OR3_X1    g038(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242_));
  INV_X1    g041(.A(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(G190gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n245_), .B(new_n241_), .C1(G183gat), .C2(G190gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G169gat), .ZN(new_n252_));
  INV_X1    g051(.A(G176gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n232_), .B1(new_n233_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n233_), .B2(new_n256_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260_));
  OAI21_X1  g059(.A(G169gat), .B1(new_n260_), .B2(KEYINPUT82), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT22), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n261_), .A2(new_n264_), .A3(new_n253_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n251_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT83), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n268_), .A3(new_n251_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n269_), .A3(new_n248_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n251_), .A2(new_n237_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n243_), .A2(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT26), .B1(new_n275_), .B2(new_n244_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n278_), .C1(KEYINPUT25), .C2(new_n243_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n246_), .B(new_n271_), .C1(new_n274_), .C2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n259_), .B1(new_n281_), .B2(new_n232_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n208_), .B1(new_n258_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n259_), .B1(new_n232_), .B2(new_n256_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n217_), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n228_), .A2(new_n229_), .B1(new_n288_), .B2(new_n220_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n226_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n231_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n214_), .A2(new_n215_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n270_), .A2(new_n291_), .A3(new_n294_), .A4(new_n280_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n284_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(new_n207_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n205_), .B1(new_n283_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n205_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n282_), .B(new_n208_), .C1(new_n232_), .C2(new_n256_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT96), .B1(new_n296_), .B2(new_n207_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n302_), .B(new_n208_), .C1(new_n284_), .C2(new_n295_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n299_), .B(new_n300_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n304_), .A3(KEYINPUT27), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n307_));
  AOI21_X1  g106(.A(new_n208_), .B1(new_n284_), .B2(new_n295_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT96), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n299_), .B1(new_n309_), .B2(new_n300_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT103), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n300_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n205_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n304_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT103), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n307_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n306_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G15gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n281_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  INV_X1    g123(.A(G43gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(new_n328_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G127gat), .B(G134gat), .Z(new_n332_));
  INV_X1    g131(.A(G120gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G113gat), .ZN(new_n334_));
  INV_X1    g133(.A(G113gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G120gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT31), .Z(new_n343_));
  NOR3_X1   g142(.A1(new_n331_), .A2(KEYINPUT86), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n329_), .A2(new_n330_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n331_), .B2(new_n343_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n346_), .A2(KEYINPUT85), .A3(new_n347_), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n344_), .A2(new_n348_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT2), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(G141gat), .A3(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT89), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n368_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n364_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n359_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n360_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(new_n365_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n357_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n353_), .B1(new_n378_), .B2(KEYINPUT1), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n356_), .A2(new_n380_), .A3(new_n357_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n342_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n364_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n385_));
  NOR4_X1   g184(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n372_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n358_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT97), .B1(new_n338_), .B2(new_n341_), .ZN(new_n390_));
  AND3_X1   g189(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT1), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n353_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n381_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n376_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n332_), .A2(new_n337_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n339_), .A2(new_n340_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n389_), .A2(new_n390_), .A3(new_n396_), .A4(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n383_), .A2(new_n384_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT99), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n383_), .A2(KEYINPUT4), .A3(new_n401_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT98), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n384_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n383_), .A2(new_n401_), .A3(KEYINPUT98), .A4(KEYINPUT4), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n383_), .A2(KEYINPUT4), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n404_), .A2(new_n411_), .A3(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(G228gat), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n374_), .A2(new_n382_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n426_), .B(new_n232_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT94), .ZN(new_n430_));
  INV_X1    g229(.A(new_n426_), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n389_), .B2(new_n396_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n289_), .A2(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n429_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n430_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n422_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n429_), .A2(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT94), .ZN(new_n440_));
  INV_X1    g239(.A(new_n422_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n429_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G22gat), .B(G50gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT28), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n389_), .A2(new_n396_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n449_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT95), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n427_), .A2(new_n447_), .A3(new_n428_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n449_), .B2(KEYINPUT29), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n445_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n444_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n438_), .A2(new_n443_), .A3(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n352_), .A2(new_n421_), .A3(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n320_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT100), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n419_), .A2(KEYINPUT33), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n404_), .A2(new_n411_), .A3(new_n466_), .A4(new_n416_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n407_), .A2(new_n384_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n383_), .A2(new_n408_), .A3(new_n401_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n417_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n315_), .A2(new_n304_), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n464_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n315_), .A2(new_n304_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT100), .A3(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n283_), .B2(new_n297_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n420_), .B(new_n478_), .C1(new_n314_), .C2(new_n477_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n461_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n459_), .A2(new_n418_), .A3(new_n419_), .A4(new_n460_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n319_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n352_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n463_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT15), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT73), .B(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT74), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G8gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT74), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n496_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n491_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n503_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n490_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT78), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n505_), .B(new_n490_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(new_n508_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G113gat), .B(G141gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G169gat), .B(G197gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n510_), .B(new_n515_), .C1(new_n511_), .C2(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT9), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G85gat), .B(G92gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n525_), .B2(KEYINPUT9), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT10), .B(G99gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(G106gat), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n535_));
  NOR2_X1   g334(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n524_), .B(KEYINPUT67), .Z(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n533_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT8), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n532_), .B1(new_n549_), .B2(new_n542_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT68), .B(G71gat), .ZN(new_n551_));
  INV_X1    g350(.A(G78gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(KEYINPUT11), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(KEYINPUT11), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n553_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n550_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n533_), .B(new_n557_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT12), .B(new_n547_), .C1(new_n558_), .C2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT12), .B1(new_n550_), .B2(KEYINPUT69), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n550_), .B2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT64), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n568_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n580_), .B2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n487_), .A2(new_n520_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n545_), .A2(new_n491_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n585_), .B(new_n591_), .C1(new_n490_), .C2(new_n545_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n590_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT72), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n594_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n600_), .B(new_n606_), .C1(new_n603_), .C2(new_n594_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n505_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n557_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT69), .B(KEYINPUT75), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n617_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n622_), .B(KEYINPUT17), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n609_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n584_), .A2(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT104), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT104), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n420_), .A2(new_n492_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n601_), .A2(new_n604_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n628_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n584_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n421_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n639_), .A3(new_n643_), .ZN(G1324gat));
  NAND4_X1  g443(.A1(new_n631_), .A2(new_n493_), .A3(new_n320_), .A4(new_n632_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n642_), .B2(new_n319_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n649_), .B(new_n651_), .ZN(G1325gat));
  OR3_X1    g451(.A1(new_n630_), .A2(G15gat), .A3(new_n486_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n642_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n352_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n655_), .B2(G15gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n461_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n654_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n659_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n663_), .A2(new_n664_), .B1(new_n630_), .B2(new_n665_), .ZN(G1327gat));
  NAND3_X1  g465(.A1(new_n582_), .A2(new_n519_), .A3(new_n628_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n478_), .B1(new_n314_), .B2(new_n477_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n474_), .A2(new_n475_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n464_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n660_), .B1(new_n672_), .B2(new_n476_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n306_), .B(new_n482_), .C1(new_n313_), .C2(new_n318_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n486_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n462_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n319_), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT43), .B(new_n608_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n480_), .A2(new_n461_), .B1(new_n319_), .B2(new_n483_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n680_), .B2(new_n352_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n681_), .B2(new_n609_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n668_), .C1(new_n678_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n487_), .B2(new_n608_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n609_), .A3(new_n679_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n667_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT109), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n668_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  INV_X1    g490(.A(new_n688_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n684_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(new_n420_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n628_), .A2(new_n640_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n584_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n420_), .A2(new_n696_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT110), .Z(new_n700_));
  OAI22_X1  g499(.A1(new_n695_), .A2(new_n696_), .B1(new_n698_), .B2(new_n700_), .ZN(G1328gat));
  NAND2_X1  g500(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n319_), .B1(new_n687_), .B2(KEYINPUT44), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n687_), .A2(KEYINPUT109), .A3(new_n688_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n691_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n319_), .A2(G36gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n584_), .A2(new_n697_), .A3(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n584_), .A2(new_n697_), .A3(new_n711_), .A4(new_n709_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n708_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n702_), .B1(new_n707_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n683_), .A2(new_n320_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n702_), .B(new_n715_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n716_), .A2(new_n721_), .ZN(G1329gat));
  XNOR2_X1  g521(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n325_), .B1(new_n698_), .B2(new_n486_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n486_), .A2(new_n325_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n730_), .B(new_n684_), .C1(new_n689_), .C2(new_n693_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n724_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n694_), .A2(new_n729_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n733_), .A2(new_n727_), .A3(new_n726_), .A4(new_n723_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1330gat));
  INV_X1    g534(.A(new_n698_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G50gat), .B1(new_n736_), .B2(new_n660_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n660_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n694_), .B2(new_n738_), .ZN(G1331gat));
  NAND3_X1  g538(.A1(new_n681_), .A2(new_n583_), .A3(new_n520_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT115), .A3(new_n641_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  INV_X1    g542(.A(new_n641_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n740_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n420_), .A2(G57gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT116), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT116), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n741_), .A2(new_n629_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n420_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n749_), .A2(new_n750_), .A3(new_n753_), .ZN(G1332gat));
  OR3_X1    g553(.A1(new_n751_), .A2(G64gat), .A3(new_n319_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n320_), .A3(new_n745_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1333gat));
  OR3_X1    g559(.A1(new_n751_), .A2(G71gat), .A3(new_n486_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n742_), .A2(new_n352_), .A3(new_n745_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT117), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1334gat));
  NAND3_X1  g569(.A1(new_n752_), .A2(new_n552_), .A3(new_n660_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n742_), .A2(new_n660_), .A3(new_n745_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G78gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G78gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(G1335gat));
  NAND2_X1  g575(.A1(new_n685_), .A2(new_n686_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n628_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n582_), .A2(new_n519_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n421_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n741_), .A2(new_n697_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n521_), .A3(new_n420_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n319_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n522_), .A3(new_n320_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n777_), .A2(new_n352_), .A3(new_n779_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G99gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n486_), .A2(new_n527_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n782_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n793_), .B(new_n794_), .Z(G1338gat));
  INV_X1    g594(.A(G106gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n782_), .A2(new_n796_), .A3(new_n660_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n777_), .A2(new_n660_), .A3(new_n779_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g602(.A1(new_n582_), .A2(new_n608_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n778_), .A2(new_n806_), .A3(new_n520_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT119), .B1(new_n628_), .B2(new_n519_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n809_));
  NAND4_X1  g608(.A1(new_n805_), .A2(new_n807_), .A3(new_n808_), .A4(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n809_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n804_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n576_), .A2(new_n519_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n576_), .B2(new_n519_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n566_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n567_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n561_), .A2(new_n563_), .A3(KEYINPUT55), .A4(new_n566_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n575_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT56), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(new_n575_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n819_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n511_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n515_), .B1(new_n829_), .B2(new_n509_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n504_), .A2(new_n507_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n509_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n518_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n577_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n828_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT122), .B(new_n815_), .C1(new_n835_), .C2(new_n640_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n640_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n576_), .B(new_n833_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n608_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n841_), .B2(new_n840_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n836_), .A2(new_n839_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n814_), .B1(new_n844_), .B2(new_n628_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n320_), .A2(new_n486_), .A3(new_n421_), .A4(new_n660_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n335_), .A3(new_n519_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n628_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n814_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT59), .A3(new_n847_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n520_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n850_), .B1(new_n857_), .B2(new_n335_), .ZN(G1340gat));
  OAI21_X1  g657(.A(new_n333_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n849_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n333_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n582_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n333_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(new_n863_), .A3(new_n778_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n628_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n849_), .A2(new_n867_), .A3(new_n640_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n608_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  NAND4_X1  g669(.A1(new_n319_), .A2(new_n486_), .A3(new_n420_), .A4(new_n660_), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(KEYINPUT124), .Z(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(new_n872_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n873_), .A2(G141gat), .A3(new_n520_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G141gat), .B1(new_n873_), .B2(new_n520_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1344gat));
  OR3_X1    g675(.A1(new_n873_), .A2(G148gat), .A3(new_n582_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G148gat), .B1(new_n873_), .B2(new_n582_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n853_), .A2(new_n778_), .A3(new_n872_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n873_), .B2(new_n608_), .ZN(new_n883_));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n640_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n873_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n845_), .A2(new_n520_), .A3(new_n319_), .A4(new_n462_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n263_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n853_), .A2(new_n519_), .A3(new_n320_), .A4(new_n676_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n252_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(G1348gat));
  NAND4_X1  g692(.A1(new_n853_), .A2(new_n583_), .A3(new_n320_), .A4(new_n676_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g694(.A1(new_n853_), .A2(new_n320_), .A3(new_n676_), .A4(new_n778_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(new_n243_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n234_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1350gat));
  NOR2_X1   g698(.A1(new_n845_), .A2(new_n319_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(new_n235_), .A3(new_n676_), .A4(new_n640_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n845_), .A2(new_n319_), .A3(new_n462_), .A4(new_n608_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n244_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n352_), .A2(new_n482_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n853_), .A2(new_n519_), .A3(new_n320_), .A4(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n900_), .A2(new_n583_), .A3(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G204gat), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n900_), .A2(new_n286_), .A3(new_n583_), .A4(new_n904_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1353gat));
  AOI21_X1  g709(.A(new_n628_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n900_), .A2(new_n904_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT126), .Z(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n900_), .A2(new_n904_), .A3(new_n911_), .A4(new_n915_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1354gat));
  AND2_X1   g718(.A1(new_n900_), .A2(new_n904_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n608_), .A2(new_n209_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n900_), .A2(new_n640_), .A3(new_n904_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n922_), .B1(new_n923_), .B2(new_n209_), .ZN(G1355gat));
endmodule


