//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT66), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(KEYINPUT66), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(new_n210_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT10), .B(G99gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(G106gat), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G85gat), .B2(G92gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(G92gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT9), .B1(new_n227_), .B2(G85gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n231_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NOR4_X1   g034(.A1(new_n232_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT69), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(new_n234_), .A3(KEYINPUT67), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT7), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n231_), .A2(new_n238_), .A3(new_n234_), .A4(KEYINPUT67), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n243_), .A3(new_n220_), .ZN(new_n244_));
  AND2_X1   g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G85gat), .A2(G92gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n217_), .A2(new_n218_), .A3(new_n210_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n210_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n240_), .B(new_n242_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n240_), .A2(new_n242_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n220_), .A3(KEYINPUT68), .ZN(new_n257_));
  INV_X1    g056(.A(new_n247_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n254_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  AOI211_X1 g059(.A(new_n209_), .B(new_n230_), .C1(new_n249_), .C2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n209_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n255_), .A2(KEYINPUT69), .B1(new_n216_), .B2(new_n219_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n258_), .B1(new_n263_), .B2(new_n243_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT8), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n259_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n256_), .B2(new_n220_), .ZN(new_n267_));
  OAI22_X1  g066(.A1(new_n264_), .A2(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n230_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n262_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT12), .B1(new_n261_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G230gat), .A2(G233gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n266_), .A2(new_n267_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n265_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n269_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n209_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n230_), .B1(new_n249_), .B2(new_n260_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n262_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n272_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291_));
  INV_X1    g090(.A(new_n289_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n279_), .A2(new_n284_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n285_), .A2(KEYINPUT70), .A3(new_n289_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n294_), .A2(new_n295_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT13), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G113gat), .B(G141gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT81), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT82), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G169gat), .B(G197gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT78), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n308_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT79), .ZN(new_n315_));
  XOR2_X1   g114(.A(G1gat), .B(G8gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G29gat), .B(G36gat), .Z(new_n318_));
  XOR2_X1   g117(.A(G43gat), .B(G50gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n316_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n315_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n315_), .A2(new_n323_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n320_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n307_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT15), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n320_), .B(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n325_), .A2(new_n331_), .A3(new_n326_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n315_), .A2(new_n323_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n321_), .B1(new_n333_), .B2(new_n324_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n307_), .B(KEYINPUT80), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OR3_X1    g135(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n306_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n306_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(new_n328_), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G169gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT83), .B(G183gat), .ZN(new_n346_));
  INV_X1    g145(.A(G190gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n345_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT84), .B1(G169gat), .B2(G176gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n355_), .A2(new_n356_), .B1(new_n364_), .B2(KEYINPUT85), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(KEYINPUT85), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n357_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n349_), .B(KEYINPUT23), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT24), .B1(new_n362_), .B2(new_n363_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT86), .B1(new_n373_), .B2(new_n351_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n352_), .B1(new_n367_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G197gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G204gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT92), .ZN(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G197gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT92), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n377_), .A3(G204gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n379_), .A2(new_n383_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT21), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n381_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT21), .ZN(new_n390_));
  XOR2_X1   g189(.A(G211gat), .B(G218gat), .Z(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(KEYINPUT21), .A3(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n376_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT19), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT97), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(KEYINPUT97), .ZN(new_n403_));
  AOI21_X1  g202(.A(G176gat), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n351_), .A2(new_n405_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n356_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n353_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n353_), .A2(KEYINPUT96), .A3(new_n408_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n407_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n369_), .A2(new_n364_), .A3(new_n371_), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n404_), .A2(new_n406_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n396_), .B(new_n400_), .C1(new_n395_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n399_), .B1(new_n415_), .B2(new_n395_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n394_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n352_), .C1(new_n367_), .C2(new_n375_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n417_), .B1(new_n422_), .B2(new_n398_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n398_), .ZN(new_n424_));
  AOI211_X1 g223(.A(KEYINPUT98), .B(new_n424_), .C1(new_n418_), .C2(new_n421_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n416_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G8gat), .B(G36gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n431_), .B(new_n416_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n376_), .B2(new_n395_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n415_), .A2(KEYINPUT101), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT101), .ZN(new_n440_));
  OAI221_X1 g239(.A(new_n440_), .B1(new_n414_), .B2(new_n413_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n441_), .A3(new_n420_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n424_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n422_), .A2(new_n398_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n436_), .B1(new_n445_), .B2(new_n432_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n435_), .A2(new_n436_), .B1(new_n446_), .B2(new_n434_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G22gat), .B(G50gat), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n450_));
  XOR2_X1   g249(.A(G155gat), .B(G162gat), .Z(new_n451_));
  INV_X1    g250(.A(KEYINPUT1), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n454_));
  INV_X1    g253(.A(G141gat), .ZN(new_n455_));
  INV_X1    g254(.A(G148gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n456_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n453_), .A2(new_n454_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT3), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n464_), .B(new_n466_), .C1(new_n457_), .C2(KEYINPUT2), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n451_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n460_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n450_), .B1(new_n469_), .B2(KEYINPUT29), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n469_), .A2(KEYINPUT29), .A3(new_n450_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n449_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n448_), .A3(new_n470_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT94), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT95), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT94), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n460_), .A2(new_n468_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n395_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT93), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(G228gat), .B1(KEYINPUT90), .B2(G233gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(KEYINPUT90), .B2(G233gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n395_), .B2(KEYINPUT89), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n395_), .B(new_n485_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n473_), .A2(new_n475_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT94), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n480_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n477_), .A2(new_n494_), .A3(new_n497_), .A4(new_n479_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G127gat), .B(G134gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G120gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n469_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n460_), .A2(new_n468_), .A3(new_n505_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT4), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n469_), .A2(new_n510_), .A3(new_n506_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n502_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G29gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G85gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT0), .B(G57gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n502_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n512_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G71gat), .B(G99gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G43gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n376_), .B(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n525_), .A2(new_n505_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n505_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(G15gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT31), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n526_), .A2(new_n533_), .A3(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n447_), .A2(new_n501_), .A3(new_n522_), .A4(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n521_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n509_), .A2(new_n502_), .A3(new_n511_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n516_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n507_), .A2(new_n517_), .A3(new_n508_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n520_), .A2(KEYINPUT33), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n516_), .C1(new_n512_), .C2(new_n518_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n434_), .A3(new_n433_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT102), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n416_), .B(new_n550_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT102), .B(new_n551_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n554_), .A2(new_n521_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n540_), .A2(new_n447_), .B1(new_n558_), .B2(new_n501_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n539_), .B1(new_n559_), .B2(new_n538_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n209_), .B(new_n561_), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n317_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n563_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(KEYINPUT17), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT74), .B1(new_n576_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n275_), .B2(new_n321_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n280_), .A2(new_n331_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT73), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n579_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n280_), .B2(new_n320_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n578_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n331_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n275_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n582_), .A2(new_n588_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n586_), .B(KEYINPUT36), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n582_), .B2(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n573_), .A2(new_n599_), .ZN(new_n600_));
  AND4_X1   g399(.A1(new_n301_), .A2(new_n343_), .A3(new_n560_), .A4(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n202_), .B1(new_n601_), .B2(new_n521_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n560_), .A2(new_n343_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n560_), .A2(KEYINPUT103), .A3(new_n343_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n580_), .A2(new_n581_), .A3(new_n578_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n591_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n596_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n582_), .A2(new_n594_), .A3(new_n588_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(KEYINPUT37), .C1(new_n611_), .C2(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT76), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n599_), .B2(new_n616_), .ZN(new_n617_));
  NOR4_X1   g416(.A1(new_n595_), .A2(new_n598_), .A3(KEYINPUT76), .A4(KEYINPUT37), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n614_), .B(KEYINPUT77), .C1(new_n617_), .C2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n572_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n607_), .A2(new_n625_), .A3(new_n301_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT104), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT104), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n627_), .A2(new_n202_), .A3(new_n521_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n602_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n630_), .B2(new_n629_), .ZN(G1324gat));
  INV_X1    g431(.A(new_n447_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n627_), .A2(new_n308_), .A3(new_n633_), .A4(new_n628_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n308_), .B1(new_n601_), .B2(new_n633_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1325gat));
  INV_X1    g442(.A(new_n626_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n530_), .A3(new_n538_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n601_), .A2(new_n538_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G15gat), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT107), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT107), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n645_), .B1(new_n651_), .B2(new_n652_), .ZN(G1326gat));
  INV_X1    g452(.A(G22gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n501_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n601_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT42), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n644_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  NAND2_X1  g458(.A1(new_n297_), .A2(new_n300_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n599_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n572_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G29gat), .B1(new_n664_), .B2(new_n521_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n621_), .A2(new_n622_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n666_), .B(new_n560_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n560_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n621_), .A2(new_n667_), .A3(new_n622_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT43), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n301_), .A2(new_n573_), .A3(new_n343_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n677_), .B(new_n674_), .C1(new_n669_), .C2(new_n672_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n521_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n665_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n679_), .B2(new_n633_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n447_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n664_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n661_), .A2(new_n663_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n686_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT45), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n682_), .B1(new_n684_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n687_), .A2(new_n690_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n676_), .A2(new_n678_), .A3(new_n447_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n693_), .B(KEYINPUT46), .C1(new_n694_), .C2(new_n683_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1329gat));
  NAND3_X1  g495(.A1(new_n661_), .A2(new_n538_), .A3(new_n663_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698_));
  INV_X1    g497(.A(G43gat), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR4_X1   g501(.A1(new_n676_), .A2(new_n678_), .A3(new_n699_), .A4(new_n537_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT47), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n679_), .A2(G43gat), .A3(new_n538_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n705_), .B(new_n706_), .C1(new_n701_), .C2(new_n700_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n664_), .B2(new_n655_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n655_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n679_), .B2(new_n710_), .ZN(G1331gat));
  AOI21_X1  g510(.A(new_n343_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n560_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n600_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n522_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n713_), .A2(new_n625_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n521_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1332gat));
  NOR2_X1   g519(.A1(new_n447_), .A2(G64gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n712_), .A2(new_n633_), .A3(new_n560_), .A4(new_n600_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G64gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT111), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n727_), .A3(G64gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n726_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n723_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n715_), .B2(new_n537_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n537_), .A2(G71gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT115), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n717_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n714_), .B2(new_n655_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT50), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n717_), .A2(new_n744_), .A3(new_n655_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1335gat));
  AND2_X1   g547(.A1(new_n713_), .A2(new_n663_), .ZN(new_n749_));
  INV_X1    g548(.A(G85gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n521_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n712_), .A2(new_n573_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n669_), .A2(new_n672_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n669_), .B2(new_n672_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n757_), .A2(new_n522_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n759_), .B2(new_n750_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT118), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n751_), .C1(new_n759_), .C2(new_n750_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1336gat));
  AOI21_X1  g563(.A(G92gat), .B1(new_n749_), .B2(new_n633_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n757_), .A2(new_n758_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n633_), .A2(new_n227_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(G1337gat));
  INV_X1    g567(.A(new_n221_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n749_), .A2(new_n769_), .A3(new_n538_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n757_), .A2(new_n537_), .A3(new_n758_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n238_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n770_), .C1(new_n771_), .C2(new_n238_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  XNOR2_X1  g575(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n754_), .A2(new_n655_), .A3(new_n673_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n713_), .A2(new_n234_), .A3(new_n655_), .A4(new_n663_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT119), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(new_n779_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n778_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(new_n780_), .A3(new_n782_), .A4(new_n777_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n625_), .A2(new_n789_), .A3(new_n301_), .A4(new_n342_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n301_), .A2(new_n342_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT54), .B1(new_n791_), .B2(new_n624_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n285_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n342_), .B1(new_n794_), .B2(new_n292_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n272_), .B1(new_n271_), .B2(new_n278_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n279_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n271_), .A2(KEYINPUT55), .A3(new_n272_), .A4(new_n278_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n289_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n802_), .B(new_n292_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n795_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n322_), .A2(new_n327_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n306_), .B1(new_n805_), .B2(new_n335_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT121), .B1(new_n332_), .B2(new_n334_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n336_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n332_), .A2(new_n334_), .A3(KEYINPUT121), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n329_), .A2(new_n337_), .A3(new_n306_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n294_), .A2(new_n812_), .A3(KEYINPUT122), .A4(new_n295_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n294_), .A2(new_n295_), .A3(new_n812_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n804_), .A2(new_n813_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n662_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT123), .B(KEYINPUT57), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(KEYINPUT57), .A3(new_n662_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n810_), .A2(new_n293_), .A3(new_n811_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT58), .B(new_n823_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(new_n621_), .A3(new_n622_), .A4(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n573_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n793_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n633_), .A2(new_n655_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n521_), .A3(new_n538_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n820_), .A2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n822_), .A2(new_n828_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n818_), .A2(KEYINPUT124), .A3(new_n819_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n573_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n833_), .B1(new_n841_), .B2(new_n793_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n343_), .B(new_n835_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G113gat), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n846_), .A3(new_n343_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1340gat));
  OAI211_X1 g647(.A(new_n660_), .B(new_n835_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n301_), .A2(KEYINPUT60), .ZN(new_n851_));
  MUX2_X1   g650(.A(new_n851_), .B(KEYINPUT60), .S(G120gat), .Z(new_n852_));
  NAND2_X1  g651(.A1(new_n842_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n842_), .B2(new_n572_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n831_), .A2(new_n834_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n842_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n572_), .A2(G127gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT125), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n855_), .B1(new_n858_), .B2(new_n860_), .ZN(G1342gat));
  OAI211_X1 g660(.A(new_n666_), .B(new_n835_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G134gat), .ZN(new_n863_));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n842_), .A2(new_n864_), .A3(new_n599_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n841_), .A2(new_n793_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n633_), .A2(new_n501_), .A3(new_n522_), .A4(new_n538_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n343_), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n660_), .A3(new_n868_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n867_), .A2(new_n572_), .A3(new_n868_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n867_), .A2(new_n876_), .A3(new_n599_), .A4(new_n868_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n867_), .A2(new_n666_), .A3(new_n868_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n876_), .ZN(G1347gat));
  NOR3_X1   g678(.A1(new_n447_), .A2(new_n521_), .A3(new_n537_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n501_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n793_), .B2(new_n830_), .ZN(new_n882_));
  AOI211_X1 g681(.A(KEYINPUT62), .B(new_n360_), .C1(new_n882_), .C2(new_n343_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n343_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(G169gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n402_), .A2(new_n403_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n882_), .A2(new_n343_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n883_), .B1(new_n886_), .B2(new_n888_), .ZN(G1348gat));
  NAND3_X1  g688(.A1(new_n660_), .A2(G176gat), .A3(new_n880_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n655_), .B(new_n890_), .C1(new_n841_), .C2(new_n793_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n881_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n831_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n361_), .B1(new_n893_), .B2(new_n301_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n361_), .C1(new_n893_), .C2(new_n301_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n891_), .B1(new_n895_), .B2(new_n897_), .ZN(G1349gat));
  NAND4_X1  g697(.A1(new_n867_), .A2(new_n572_), .A3(new_n501_), .A4(new_n880_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n572_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n899_), .A2(new_n346_), .B1(new_n882_), .B2(new_n900_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n893_), .B2(new_n623_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n882_), .A2(new_n599_), .A3(new_n356_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n633_), .A2(new_n540_), .A3(new_n537_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n841_), .B2(new_n793_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n343_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n660_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n911_));
  INV_X1    g710(.A(G211gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(KEYINPUT127), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n913_), .B(new_n573_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n906_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT127), .B1(new_n911_), .B2(new_n912_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1354gat));
  INV_X1    g716(.A(new_n906_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G218gat), .B1(new_n918_), .B2(new_n623_), .ZN(new_n919_));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n906_), .A2(new_n920_), .A3(new_n599_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1355gat));
endmodule


