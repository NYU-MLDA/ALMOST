//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  INV_X1    g001(.A(G230gat), .ZN(new_n203_));
  INV_X1    g002(.A(G233gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206_));
  AND2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT67), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n212_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  OAI22_X1  g025(.A1(new_n226_), .A2(KEYINPUT69), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n222_), .A2(KEYINPUT7), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n225_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n211_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n213_), .A2(new_n214_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT70), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n225_), .B(new_n232_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n224_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n222_), .A2(KEYINPUT7), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(KEYINPUT69), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n232_), .B1(new_n238_), .B2(new_n225_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n231_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n209_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n230_), .B1(new_n241_), .B2(KEYINPUT8), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT9), .B1(new_n207_), .B2(new_n208_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT66), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n207_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(new_n215_), .A3(new_n220_), .A4(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT65), .B(G106gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT10), .B(G99gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT64), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(new_n249_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n250_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT64), .B1(new_n254_), .B2(new_n255_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n243_), .A2(new_n246_), .B1(new_n207_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(new_n221_), .A3(new_n264_), .A4(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n206_), .B1(new_n242_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n231_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n229_), .A2(KEYINPUT70), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n233_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n209_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT8), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n230_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n258_), .A2(new_n266_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT71), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n268_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n281_));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT72), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT73), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n268_), .A2(new_n286_), .A3(new_n277_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n268_), .B2(new_n277_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n205_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n275_), .A2(new_n276_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n285_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT12), .A3(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n290_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n205_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G120gat), .B(G148gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT5), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  OAI21_X1  g106(.A(new_n202_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n294_), .A2(new_n302_), .A3(KEYINPUT74), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n314_));
  NAND2_X1  g113(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(KEYINPUT75), .A3(KEYINPUT13), .A4(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G29gat), .B(G36gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G43gat), .B(G50gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G15gat), .B(G22gat), .ZN(new_n326_));
  INV_X1    g125(.A(G1gat), .ZN(new_n327_));
  INV_X1    g126(.A(G8gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G8gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n325_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT82), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G229gat), .A3(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n325_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(new_n332_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n325_), .B(KEYINPUT15), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n332_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT83), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G169gat), .B(G197gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n320_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n336_), .A2(new_n343_), .A3(KEYINPUT85), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n336_), .A2(KEYINPUT84), .A3(new_n343_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT84), .B1(new_n336_), .B2(new_n343_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n319_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT108), .ZN(new_n357_));
  INV_X1    g156(.A(new_n355_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n318_), .A2(KEYINPUT108), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G141gat), .B(G148gat), .Z(new_n361_));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT92), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364_));
  AND2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(KEYINPUT93), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(KEYINPUT1), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT93), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n363_), .A2(new_n367_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(KEYINPUT94), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(KEYINPUT94), .A2(KEYINPUT3), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT2), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n375_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n383_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n372_), .A2(new_n381_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n384_), .B(KEYINPUT90), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n385_), .B(KEYINPUT89), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n381_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n369_), .A2(new_n370_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(new_n366_), .C1(KEYINPUT1), .C2(new_n367_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n394_), .B2(new_n361_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n387_), .B(new_n388_), .C1(new_n391_), .C2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT101), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n372_), .A2(new_n381_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(KEYINPUT101), .A3(new_n387_), .A4(new_n388_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n388_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n404_), .B(new_n405_), .C1(KEYINPUT4), .C2(new_n401_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT0), .ZN(new_n408_));
  INV_X1    g207(.A(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n403_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT102), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n403_), .A2(new_n406_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n412_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT102), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n403_), .A2(new_n406_), .A3(new_n413_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n391_), .B(KEYINPUT31), .Z(new_n425_));
  INV_X1    g224(.A(G183gat), .ZN(new_n426_));
  INV_X1    g225(.A(G190gat), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT23), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT23), .B1(new_n426_), .B2(new_n427_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(KEYINPUT87), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(KEYINPUT87), .B2(new_n429_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G169gat), .ZN(new_n436_));
  INV_X1    g235(.A(G176gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(new_n428_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT24), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OR3_X1    g243(.A1(new_n435_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT25), .B(G183gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT86), .B1(new_n427_), .B2(KEYINPUT26), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(G190gat), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n446_), .B(new_n447_), .C1(new_n448_), .C2(KEYINPUT86), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n441_), .A2(new_n444_), .A3(new_n445_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n439_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT30), .Z(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(G15gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT88), .B(G43gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n452_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n425_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n459_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT91), .A3(new_n425_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n424_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT106), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT104), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G8gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT18), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(KEYINPUT103), .Z(new_n473_));
  XNOR2_X1  g272(.A(G197gat), .B(G204gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G211gat), .B(G218gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT21), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G204gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G197gat), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n480_), .B2(KEYINPUT95), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(new_n474_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n475_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT96), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n483_), .A2(KEYINPUT96), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n478_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n431_), .A2(new_n444_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT98), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT98), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n431_), .A2(new_n490_), .A3(new_n444_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n448_), .A2(new_n446_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n445_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n489_), .A2(KEYINPUT99), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n441_), .A2(new_n433_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n438_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n491_), .A2(new_n493_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT99), .B1(new_n498_), .B2(new_n489_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n487_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT19), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n483_), .A2(KEYINPUT96), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n477_), .B1(new_n505_), .B2(new_n484_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n451_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n500_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n504_), .B1(new_n487_), .B2(new_n451_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n498_), .A2(new_n489_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n511_), .A3(new_n496_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n503_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n468_), .B(new_n473_), .C1(new_n509_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n500_), .A2(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n502_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n491_), .A2(new_n493_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n490_), .B1(new_n431_), .B2(new_n444_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n506_), .A2(new_n520_), .A3(new_n494_), .A4(new_n496_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI211_X1 g322(.A(new_n504_), .B(new_n502_), .C1(new_n487_), .C2(new_n451_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n494_), .A2(new_n496_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n525_), .A2(KEYINPUT100), .A3(new_n506_), .A4(new_n520_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n516_), .A2(new_n527_), .A3(new_n472_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n506_), .A2(new_n511_), .A3(new_n496_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT20), .B1(new_n506_), .B2(new_n507_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n502_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n502_), .B2(new_n515_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n468_), .B1(new_n533_), .B2(new_n473_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT27), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n516_), .A2(new_n527_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n472_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT27), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n528_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G78gat), .B(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n543_));
  INV_X1    g342(.A(G228gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n204_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n487_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n543_), .B2(new_n487_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n542_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n543_), .A2(new_n487_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n545_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(new_n487_), .A3(new_n546_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT28), .B1(new_n399_), .B2(KEYINPUT29), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n395_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G22gat), .B(G50gat), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n555_), .A2(new_n557_), .A3(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n565_), .A2(new_n566_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n554_), .B(new_n549_), .C1(new_n569_), .C2(new_n556_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n467_), .B1(new_n541_), .B2(new_n572_), .ZN(new_n573_));
  AOI211_X1 g372(.A(KEYINPUT106), .B(new_n571_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n466_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT107), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n416_), .A2(new_n422_), .B1(new_n570_), .B2(new_n568_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n541_), .A2(KEYINPUT105), .A3(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n472_), .A2(KEYINPUT32), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n533_), .A2(new_n580_), .ZN(new_n581_));
  OAI221_X1 g380(.A(new_n581_), .B1(new_n536_), .B2(new_n580_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n538_), .A2(new_n528_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n421_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n403_), .A2(new_n406_), .A3(KEYINPUT33), .A4(new_n413_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n401_), .A2(new_n387_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n404_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n388_), .B1(new_n401_), .B2(KEYINPUT4), .ZN(new_n589_));
  OAI221_X1 g388(.A(new_n412_), .B1(new_n587_), .B2(new_n388_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(new_n586_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n582_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n572_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n579_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT105), .B1(new_n541_), .B2(new_n578_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n465_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT107), .B(new_n466_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n577_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT36), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT77), .B(KEYINPUT34), .Z(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n278_), .A2(KEYINPUT79), .A3(new_n337_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT79), .B1(new_n278_), .B2(new_n337_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n607_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT80), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n339_), .B2(new_n297_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n609_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n609_), .A3(new_n616_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n603_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n601_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n621_), .A2(new_n617_), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT16), .ZN(new_n628_));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n332_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n632_), .B1(new_n287_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n287_), .B2(new_n635_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n631_), .B(new_n630_), .C1(new_n634_), .C2(new_n298_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n298_), .B2(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n626_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n360_), .A2(new_n598_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n424_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n620_), .B2(new_n625_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n602_), .B1(new_n621_), .B2(new_n617_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n623_), .A3(new_n619_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n640_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT81), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n358_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n318_), .A2(KEYINPUT76), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n318_), .A2(KEYINPUT76), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n598_), .A3(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n643_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n644_), .B1(new_n662_), .B2(new_n663_), .ZN(G1324gat));
  OAI21_X1  g463(.A(G8gat), .B1(new_n642_), .B2(new_n541_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(new_n541_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n328_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n666_), .A2(new_n667_), .B1(new_n659_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI221_X1 g471(.A(KEYINPUT40), .B1(new_n659_), .B2(new_n669_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n642_), .B2(new_n465_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n659_), .A2(G15gat), .A3(new_n465_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(G1326gat));
  OAI21_X1  g479(.A(G22gat), .B1(new_n642_), .B2(new_n572_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT42), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n572_), .A2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n659_), .B2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n626_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n652_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n319_), .A2(new_n355_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n595_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n579_), .A3(new_n593_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n689_), .A2(new_n465_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n687_), .B1(new_n690_), .B2(new_n597_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n692_), .A2(G29gat), .A3(new_n643_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n652_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n598_), .A2(new_n695_), .A3(new_n650_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n598_), .B2(new_n650_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n694_), .B(KEYINPUT44), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n424_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G29gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n693_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n700_), .A2(new_n668_), .A3(new_n701_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n541_), .A2(G36gat), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n691_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n691_), .B2(new_n714_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n709_), .B1(new_n711_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n717_), .B(new_n708_), .C1(new_n710_), .C2(G36gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(new_n465_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n700_), .A2(G43gat), .A3(new_n722_), .A4(new_n701_), .ZN(new_n723_));
  INV_X1    g522(.A(G43gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n692_), .B2(new_n465_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n691_), .B2(new_n571_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n701_), .A2(G50gat), .A3(new_n571_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n700_), .ZN(G1331gat));
  AOI21_X1  g529(.A(new_n355_), .B1(new_n690_), .B2(new_n597_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n654_), .A2(new_n319_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n409_), .A3(new_n424_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n658_), .A2(new_n640_), .A3(new_n626_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n731_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n643_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n737_), .B2(new_n541_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n734_), .A2(new_n743_), .A3(new_n668_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n737_), .B2(new_n465_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n734_), .A2(new_n748_), .A3(new_n722_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n572_), .A2(G78gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT114), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n732_), .A2(new_n733_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n736_), .A2(new_n571_), .A3(new_n731_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT115), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n753_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n658_), .A2(new_n652_), .A3(new_n685_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n732_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n411_), .A3(new_n424_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n319_), .A2(new_n355_), .A3(new_n652_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT116), .B(new_n766_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n643_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n411_), .B2(new_n771_), .ZN(G1336gat));
  INV_X1    g571(.A(G92gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n764_), .A2(new_n773_), .A3(new_n668_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n541_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(new_n775_), .ZN(G1337gat));
  AOI21_X1  g575(.A(new_n465_), .B1(new_n256_), .B2(new_n253_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n732_), .A2(new_n763_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n465_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n223_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n778_), .C1(new_n779_), .C2(new_n223_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1338gat));
  NAND4_X1  g583(.A1(new_n732_), .A2(new_n259_), .A3(new_n571_), .A4(new_n763_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n571_), .B(new_n766_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G106gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G106gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n785_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT12), .B1(new_n278_), .B2(new_n287_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n290_), .A2(new_n299_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n205_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n290_), .B(new_n299_), .C1(new_n291_), .C2(KEYINPUT12), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT117), .A3(new_n205_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT55), .B1(new_n801_), .B2(new_n205_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n296_), .A2(new_n300_), .A3(new_n805_), .A4(new_n301_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n307_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n810_), .B(new_n309_), .C1(new_n803_), .C2(new_n807_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n311_), .B(new_n355_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n800_), .A2(new_n802_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n815_), .B2(new_n309_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n307_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(KEYINPUT118), .A3(new_n311_), .A4(new_n355_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n335_), .A2(new_n342_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n342_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n349_), .B1(new_n340_), .B2(new_n821_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n348_), .A2(new_n350_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n313_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n819_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n685_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT119), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n818_), .A2(new_n311_), .A3(new_n823_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n650_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n816_), .A2(new_n817_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n831_), .B2(new_n823_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT57), .B1(new_n825_), .B2(new_n685_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n640_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n650_), .A2(new_n355_), .A3(new_n640_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n319_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(new_n319_), .A3(KEYINPUT54), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n424_), .B(new_n722_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n848_), .B(new_n845_), .C1(new_n836_), .C2(new_n843_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n795_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n830_), .A2(new_n832_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n812_), .A2(new_n813_), .B1(new_n313_), .B2(new_n823_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n626_), .B1(new_n852_), .B2(new_n819_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n825_), .A2(new_n685_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n652_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n846_), .B1(new_n858_), .B2(new_n842_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n848_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n846_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT120), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n358_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n850_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n859_), .B2(new_n358_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1340gat));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n868_));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n318_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n844_), .A2(new_n846_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n658_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n869_), .ZN(G1341gat));
  NAND2_X1  g673(.A1(new_n652_), .A2(G127gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT121), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n850_), .A2(new_n862_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n859_), .B2(new_n640_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1342gat));
  XOR2_X1   g679(.A(KEYINPUT122), .B(G134gat), .Z(new_n881_));
  NOR2_X1   g680(.A1(new_n651_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n850_), .A2(new_n862_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n859_), .B2(new_n685_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n858_), .A2(new_n842_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n424_), .A2(new_n571_), .A3(new_n465_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n887_), .A2(new_n668_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n355_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g690(.A(new_n658_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(G148gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n652_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(G162gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n889_), .A2(new_n899_), .A3(new_n626_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n889_), .A2(new_n650_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1347gat));
  INV_X1    g701(.A(new_n466_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n903_), .A2(new_n541_), .A3(new_n571_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n887_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n355_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G169gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n907_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n906_), .A2(new_n355_), .A3(new_n436_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n844_), .A2(new_n318_), .A3(new_n904_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n437_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(KEYINPUT124), .A3(new_n437_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n658_), .A2(new_n437_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n917_), .A2(new_n918_), .B1(new_n906_), .B2(new_n919_), .ZN(G1349gat));
  NAND2_X1  g719(.A1(new_n906_), .A2(new_n652_), .ZN(new_n921_));
  MUX2_X1   g720(.A(new_n446_), .B(G183gat), .S(new_n921_), .Z(G1350gat));
  NAND2_X1  g721(.A1(new_n626_), .A2(new_n448_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT125), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n906_), .A2(new_n924_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n887_), .A2(new_n651_), .A3(new_n905_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n427_), .B2(new_n926_), .ZN(G1351gat));
  NAND3_X1  g726(.A1(new_n668_), .A2(new_n465_), .A3(new_n578_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n355_), .B(new_n929_), .C1(new_n858_), .C2(new_n842_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT127), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n928_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n933_), .A2(KEYINPUT126), .A3(new_n934_), .A4(new_n355_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(KEYINPUT126), .B1(new_n933_), .B2(new_n355_), .ZN(new_n937_));
  INV_X1    g736(.A(G197gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n936_), .A2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n932_), .B(new_n935_), .C1(new_n938_), .C2(new_n937_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n933_), .A2(new_n892_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g743(.A(new_n933_), .ZN(new_n945_));
  OAI22_X1  g744(.A1(new_n945_), .A2(new_n640_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT63), .B(G211gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n933_), .A2(new_n652_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n945_), .B2(new_n651_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n685_), .A2(G218gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n945_), .B2(new_n951_), .ZN(G1355gat));
endmodule


