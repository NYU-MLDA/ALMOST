//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT73), .B(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT22), .B1(new_n207_), .B2(KEYINPUT72), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G169gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n206_), .B(new_n208_), .C1(KEYINPUT72), .C2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(G183gat), .C2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT25), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G190gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n233_), .A2(new_n234_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n227_), .B(new_n232_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n228_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT71), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n218_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT21), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n245_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n244_), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n245_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n248_), .A2(new_n251_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255_));
  INV_X1    g054(.A(KEYINPUT83), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(KEYINPUT83), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  AOI211_X1 g060(.A(new_n203_), .B(new_n205_), .C1(new_n243_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT22), .B(G169gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n206_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n267_), .A2(new_n268_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT85), .B1(new_n269_), .B2(new_n235_), .ZN(new_n270_));
  AND4_X1   g069(.A1(KEYINPUT85), .A2(new_n235_), .A3(new_n227_), .A4(new_n232_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n272_), .B2(new_n261_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n266_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n235_), .A2(new_n227_), .A3(new_n232_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(KEYINPUT85), .A3(new_n235_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n261_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT87), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n262_), .A2(new_n273_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n262_), .A2(new_n273_), .A3(KEYINPUT88), .A4(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n241_), .A2(KEYINPUT71), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n235_), .A2(new_n236_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n269_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n289_), .A2(new_n260_), .A3(new_n254_), .A4(new_n218_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n290_), .B(KEYINPUT20), .C1(new_n279_), .C2(new_n280_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n205_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(KEYINPUT86), .A3(new_n205_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  NAND3_X1  g099(.A1(new_n286_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(G141gat), .ZN(new_n312_));
  INV_X1    g111(.A(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  AND4_X1   g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n309_), .A2(new_n323_), .A3(new_n305_), .ZN(new_n324_));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT76), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n315_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT81), .A3(new_n261_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT80), .ZN(new_n332_));
  INV_X1    g131(.A(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(new_n336_), .A3(new_n261_), .A4(KEYINPUT81), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT78), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT77), .B(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n342_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n344_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n319_), .A2(new_n317_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n315_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n341_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n350_), .B1(new_n341_), .B2(new_n355_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n341_), .A2(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n363_), .B2(new_n356_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n338_), .B(new_n340_), .C1(new_n360_), .C2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT84), .B(new_n359_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n359_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n367_), .A3(new_n356_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n338_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n366_), .B(new_n368_), .C1(new_n369_), .C2(new_n339_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n243_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT20), .B1(new_n372_), .B2(new_n280_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n280_), .A2(new_n266_), .A3(new_n275_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n205_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n205_), .B2(new_n291_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n300_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n202_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n301_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G134gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G127gat), .ZN(new_n381_));
  INV_X1    g180(.A(G127gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G134gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G120gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G113gat), .ZN(new_n386_));
  INV_X1    g185(.A(G113gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G120gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n381_), .A2(new_n383_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n390_), .A2(KEYINPUT74), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT74), .B1(new_n390_), .B2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n394_), .B(KEYINPUT31), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G15gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT30), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  INV_X1    g202(.A(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n402_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(new_n372_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n397_), .A2(new_n398_), .A3(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n390_), .A2(KEYINPUT74), .A3(new_n391_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT74), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n384_), .A2(new_n389_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n381_), .A2(new_n383_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n329_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n352_), .B(new_n315_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n415_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT4), .B1(new_n394_), .B2(new_n329_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n414_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT4), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n421_), .A2(new_n415_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n414_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n410_), .A2(new_n437_), .ZN(new_n438_));
  AND4_X1   g237(.A1(new_n304_), .A2(new_n371_), .A3(new_n379_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n286_), .A2(new_n296_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n377_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n423_), .A2(new_n424_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n427_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n434_), .B1(new_n430_), .B2(new_n425_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n428_), .B1(new_n442_), .B2(new_n427_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT33), .B1(new_n446_), .B2(new_n434_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n414_), .C1(new_n426_), .C2(new_n428_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n450_), .A3(new_n301_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n376_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n437_), .B(new_n453_), .C1(new_n440_), .C2(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n371_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n437_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n304_), .A2(new_n457_), .A3(new_n379_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT27), .B1(new_n441_), .B2(new_n301_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n379_), .A2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT89), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n439_), .B1(new_n463_), .B2(new_n410_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G29gat), .B(G36gat), .Z(new_n465_));
  XOR2_X1   g264(.A(G43gat), .B(G50gat), .Z(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT15), .Z(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n468_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n467_), .A2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n467_), .B(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G141gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G169gat), .B(G197gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n483_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G176gat), .B(G204gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G230gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT6), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  OR3_X1    g296(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G85gat), .B(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT64), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n499_), .A2(new_n507_), .A3(new_n502_), .A4(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT9), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n510_), .A2(new_n513_), .A3(new_n496_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  XOR2_X1   g319(.A(G71gat), .B(G78gat), .Z(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n494_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n517_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n509_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n506_), .A2(KEYINPUT66), .A3(new_n508_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n525_), .A2(KEYINPUT12), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n526_), .B1(new_n539_), .B2(new_n528_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n493_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n492_), .B1(new_n531_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(new_n541_), .A3(new_n492_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n543_), .B(new_n544_), .C1(KEYINPUT67), .C2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n547_));
  INV_X1    g346(.A(new_n544_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n542_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n532_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n467_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n552_), .A2(new_n553_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n468_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n536_), .B2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n554_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n558_), .C1(new_n536_), .C2(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT36), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n571_), .A3(new_n564_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n551_), .B1(new_n573_), .B2(KEYINPUT69), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n475_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n525_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n577_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n583_), .B2(new_n577_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT69), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n570_), .A2(new_n591_), .A3(KEYINPUT37), .A4(new_n572_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n574_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n464_), .A2(new_n487_), .A3(new_n550_), .A4(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT90), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n470_), .A3(new_n437_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT92), .ZN(new_n599_));
  INV_X1    g398(.A(new_n573_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n464_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n546_), .A2(new_n549_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n487_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n590_), .A3(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT93), .Z(new_n607_));
  AOI21_X1  g406(.A(new_n470_), .B1(new_n607_), .B2(new_n437_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT94), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n596_), .A2(new_n597_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT95), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n609_), .A3(new_n611_), .ZN(G1324gat));
  AND2_X1   g411(.A1(new_n304_), .A2(new_n379_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT39), .ZN(new_n615_));
  INV_X1    g414(.A(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n595_), .A2(new_n471_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g418(.A(new_n410_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n400_), .B1(new_n607_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT41), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n595_), .A2(new_n400_), .A3(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n371_), .B(KEYINPUT96), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n595_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n607_), .B2(new_n626_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT97), .B(KEYINPUT42), .Z(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT98), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n634_), .B(new_n627_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1327gat));
  NOR2_X1   g435(.A1(new_n464_), .A2(new_n487_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n590_), .A2(new_n573_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n602_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(G29gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n437_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n574_), .A2(new_n592_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n463_), .A2(new_n410_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n439_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n464_), .A2(KEYINPUT99), .A3(KEYINPUT43), .A4(new_n649_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n651_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n649_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n654_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n604_), .A2(new_n590_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n647_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n653_), .A3(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT99), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n464_), .A2(KEYINPUT43), .A3(new_n649_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n648_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n464_), .B2(new_n649_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n660_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n437_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n645_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT103), .B(new_n645_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1328gat));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n616_), .A3(new_n669_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G36gat), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n613_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n641_), .A2(new_n642_), .A3(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT104), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1329gat));
  AOI21_X1  g485(.A(G43gat), .B1(new_n643_), .B2(new_n620_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n662_), .A2(new_n669_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n410_), .A2(new_n404_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n643_), .B2(new_n626_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n371_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n688_), .B2(new_n694_), .ZN(G1331gat));
  NOR4_X1   g494(.A1(new_n464_), .A2(new_n603_), .A3(new_n602_), .A4(new_n593_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n437_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n550_), .A2(new_n487_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n590_), .ZN(new_n700_));
  NOR4_X1   g499(.A1(new_n464_), .A2(new_n699_), .A3(new_n600_), .A4(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n437_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n702_), .B2(new_n697_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n701_), .B2(new_n616_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n704_), .A3(new_n616_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n701_), .B2(new_n620_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(KEYINPUT49), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n709_), .A3(new_n620_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT106), .Z(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n701_), .B2(new_n626_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n696_), .A2(new_n716_), .A3(new_n626_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT107), .Z(G1335gat));
  NOR2_X1   g520(.A1(new_n699_), .A2(new_n590_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n668_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(new_n437_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n656_), .A2(new_n487_), .A3(new_n550_), .A4(new_n638_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n514_), .A3(new_n437_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1336gat));
  OAI21_X1  g528(.A(G92gat), .B1(new_n724_), .B2(new_n613_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n515_), .A3(new_n616_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n724_), .B2(new_n410_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n620_), .A2(new_n511_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT109), .B1(new_n727_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n727_), .A2(new_n512_), .A3(new_n693_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n667_), .B1(new_n665_), .B2(new_n648_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n693_), .B(new_n722_), .C1(new_n742_), .C2(new_n655_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n668_), .A2(KEYINPUT110), .A3(new_n693_), .A4(new_n722_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n512_), .B1(KEYINPUT111), .B2(KEYINPUT52), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n747_), .A2(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n750_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n748_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n752_), .B(new_n753_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n741_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n741_), .C1(new_n751_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n538_), .A2(new_n540_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n494_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n541_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n761_), .A2(new_n760_), .A3(new_n494_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n491_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT56), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n491_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n767_), .A2(new_n603_), .A3(new_n544_), .A4(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n486_), .B1(new_n480_), .B2(new_n478_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n476_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n479_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(KEYINPUT115), .A3(new_n773_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n776_), .A2(KEYINPUT116), .A3(new_n777_), .A4(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n770_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n573_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n548_), .B1(new_n766_), .B2(KEYINPUT56), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n783_), .A3(new_n769_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n790_), .A2(KEYINPUT58), .A3(new_n783_), .A4(new_n769_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n657_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n600_), .B1(new_n770_), .B2(new_n784_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT57), .B1(new_n796_), .B2(KEYINPUT117), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n789_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n550_), .A2(new_n593_), .A3(new_n603_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n649_), .A2(new_n590_), .A3(new_n487_), .A4(new_n602_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(KEYINPUT54), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n802_), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n798_), .A2(new_n700_), .B1(new_n805_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n616_), .A2(new_n693_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n437_), .A3(new_n620_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813_), .B2(new_n603_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n798_), .A2(new_n700_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n805_), .A2(new_n809_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n812_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(KEYINPUT59), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n603_), .A2(G113gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT118), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n822_), .B2(new_n824_), .ZN(G1340gat));
  AOI21_X1  g624(.A(new_n602_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n385_), .B1(new_n602_), .B2(KEYINPUT60), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT119), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(G120gat), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n813_), .A2(KEYINPUT120), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT120), .B1(new_n813_), .B2(new_n830_), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n826_), .A2(new_n385_), .B1(new_n831_), .B2(new_n832_), .ZN(G1341gat));
  NAND3_X1  g632(.A1(new_n813_), .A2(new_n382_), .A3(new_n590_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n700_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n382_), .ZN(G1342gat));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n380_), .B1(new_n822_), .B2(new_n657_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n813_), .A2(new_n380_), .A3(new_n600_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n649_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT121), .B(new_n839_), .C1(new_n842_), .C2(new_n380_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1343gat));
  NAND2_X1  g643(.A1(new_n693_), .A2(new_n410_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n616_), .A2(new_n725_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n817_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n487_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n312_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n602_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n313_), .ZN(G1345gat));
  OR3_X1    g650(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n700_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n700_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1346gat));
  INV_X1    g656(.A(G162gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n847_), .A2(new_n858_), .A3(new_n649_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n847_), .B2(new_n573_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n861_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n616_), .A2(new_n438_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n810_), .A2(new_n626_), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n264_), .A3(new_n603_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n626_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n817_), .A2(new_n603_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT62), .B1(new_n870_), .B2(G169gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n865_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .A3(new_n868_), .A4(new_n871_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1348gat));
  NAND2_X1  g676(.A1(new_n867_), .A2(new_n550_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n810_), .A2(new_n693_), .ZN(new_n879_));
  INV_X1    g678(.A(G176gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n866_), .A2(new_n880_), .A3(new_n602_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n878_), .A2(new_n206_), .B1(new_n879_), .B2(new_n881_), .ZN(G1349gat));
  INV_X1    g681(.A(new_n867_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n267_), .A3(new_n700_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n879_), .A2(new_n616_), .A3(new_n438_), .A4(new_n590_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n219_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n883_), .B2(new_n649_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n867_), .A2(new_n268_), .A3(new_n600_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n613_), .A2(new_n437_), .A3(new_n845_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n817_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(G197gat), .ZN(new_n892_));
  OAI22_X1  g691(.A1(new_n891_), .A2(new_n487_), .B1(KEYINPUT125), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT126), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(new_n895_), .ZN(G1352gat));
  INV_X1    g695(.A(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n550_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT127), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n897_), .A2(new_n590_), .A3(new_n901_), .A4(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n900_), .A2(KEYINPUT127), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1354gat));
  OR3_X1    g704(.A1(new_n891_), .A2(G218gat), .A3(new_n573_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G218gat), .B1(new_n891_), .B2(new_n649_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1355gat));
endmodule


