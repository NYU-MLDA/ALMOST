//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(KEYINPUT77), .A2(G1gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT77), .A2(G1gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT78), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n212_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT77), .A2(G1gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(G8gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT14), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G15gat), .B(G22gat), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n209_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n209_), .ZN(new_n225_));
  AOI211_X1 g024(.A(new_n222_), .B(new_n225_), .C1(new_n215_), .C2(new_n220_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n208_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n213_), .A2(KEYINPUT78), .A3(new_n214_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n219_), .B1(new_n218_), .B2(KEYINPUT14), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n223_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n225_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n208_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n221_), .A2(new_n223_), .A3(new_n209_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT79), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(new_n234_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239_));
  INV_X1    g038(.A(new_n236_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n236_), .B(KEYINPUT80), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n233_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n204_), .A2(KEYINPUT15), .A3(new_n207_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT15), .B1(new_n204_), .B2(new_n207_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n227_), .B(new_n243_), .C1(new_n244_), .C2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G169gat), .B(G197gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  NAND4_X1  g050(.A1(new_n242_), .A2(KEYINPUT82), .A3(new_n248_), .A4(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n239_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT79), .B(new_n236_), .C1(new_n227_), .C2(new_n234_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n248_), .B(new_n251_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n242_), .A2(new_n248_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n251_), .B(KEYINPUT81), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(G71gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G99gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT85), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n266_), .B(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G183gat), .A3(G190gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT23), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n271_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT25), .B(G183gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT83), .B1(new_n283_), .B2(G190gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n282_), .B(new_n284_), .C1(new_n285_), .C2(KEYINPUT83), .ZN(new_n286_));
  NOR3_X1   g085(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT24), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n286_), .B(new_n288_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n281_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT30), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT86), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(KEYINPUT86), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n269_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n297_), .B2(new_n269_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT87), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT87), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT88), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT31), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n300_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n300_), .A2(new_n312_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT101), .ZN(new_n318_));
  XOR2_X1   g117(.A(G64gat), .B(G92gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(G204gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G197gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT21), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(KEYINPUT93), .B2(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n323_), .B2(G204gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n327_), .B(new_n328_), .C1(new_n332_), .C2(KEYINPUT21), .ZN(new_n333_));
  INV_X1    g132(.A(new_n328_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(KEYINPUT21), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n294_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n289_), .A2(new_n290_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G169gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT96), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n340_), .B2(new_n290_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n280_), .B1(new_n277_), .B2(new_n273_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT97), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n287_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n345_), .A2(new_n275_), .A3(new_n278_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n292_), .B1(new_n291_), .B2(KEYINPUT95), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(KEYINPUT95), .B2(new_n291_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n337_), .B(KEYINPUT20), .C1(new_n350_), .C2(new_n336_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n336_), .B2(new_n294_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n350_), .A2(new_n358_), .A3(new_n336_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n341_), .A2(new_n343_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n333_), .A2(new_n335_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT98), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n357_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(new_n354_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT99), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n356_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT99), .B1(new_n363_), .B2(new_n354_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n322_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n358_), .B1(new_n350_), .B2(new_n336_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT98), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n365_), .B(new_n355_), .C1(new_n371_), .C2(new_n357_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n356_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n322_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n316_), .B1(new_n368_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n366_), .A2(new_n322_), .A3(new_n367_), .ZN(new_n378_));
  MUX2_X1   g177(.A(new_n351_), .B(new_n363_), .S(new_n354_), .Z(new_n379_));
  AOI21_X1  g178(.A(new_n316_), .B1(new_n379_), .B2(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT90), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(G155gat), .B2(G162gat), .ZN(new_n384_));
  OR3_X1    g183(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT2), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  OR3_X1    g191(.A1(KEYINPUT89), .A2(G141gat), .A3(G148gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n393_), .A2(new_n394_), .B1(G141gat), .B2(G148gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT1), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n383_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n309_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n392_), .A2(new_n307_), .A3(new_n308_), .A4(new_n398_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(KEYINPUT4), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT102), .Z(new_n404_));
  OAI211_X1 g203(.A(new_n402_), .B(new_n404_), .C1(KEYINPUT4), .C2(new_n400_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n400_), .A2(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT0), .B(G57gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n405_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT92), .A3(new_n336_), .ZN(new_n418_));
  AND2_X1   g217(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(G233gat), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G78gat), .ZN(new_n422_));
  INV_X1    g221(.A(G106gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n418_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G22gat), .B(G50gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n428_), .A2(new_n429_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n427_), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n426_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n426_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n416_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n377_), .A2(new_n381_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n374_), .A2(new_n375_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n415_), .A2(KEYINPUT33), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n405_), .A2(new_n407_), .A3(new_n443_), .A4(new_n412_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n402_), .B(new_n403_), .C1(KEYINPUT4), .C2(new_n400_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n412_), .B1(new_n406_), .B2(new_n404_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n442_), .A2(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n378_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n379_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n450_), .B(new_n416_), .C1(new_n374_), .C2(new_n449_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n440_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n439_), .B1(new_n452_), .B2(KEYINPUT103), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT103), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n454_), .B(new_n440_), .C1(new_n448_), .C2(new_n451_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n315_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n377_), .A2(new_n381_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n315_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n416_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n440_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n262_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G57gat), .B(G64gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT69), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(KEYINPUT66), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT66), .ZN(new_n479_));
  AND2_X1   g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n476_), .A2(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT66), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT10), .B(G99gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(G106gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n474_), .B1(new_n485_), .B2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(G85gat), .B(G92gat), .C1(new_n482_), .C2(KEYINPUT9), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n482_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n483_), .ZN(new_n497_));
  AND2_X1   g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n500_), .A2(new_n423_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(KEYINPUT67), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G85gat), .B(G92gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT8), .B(new_n504_), .C1(new_n508_), .C2(new_n490_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  OR3_X1    g309(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n488_), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n511_), .B(new_n505_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n504_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n471_), .B(new_n473_), .C1(new_n503_), .C2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n497_), .A2(new_n501_), .A3(KEYINPUT67), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT67), .B1(new_n497_), .B2(new_n501_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT8), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n470_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n518_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n525_), .A2(new_n502_), .A3(new_n493_), .A4(new_n470_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n463_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n471_), .B1(new_n503_), .B2(new_n517_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n521_), .A2(KEYINPUT68), .A3(new_n525_), .A4(new_n470_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n529_), .A2(new_n532_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n527_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT70), .A4(new_n518_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n546_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT13), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT34), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT74), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n559_), .B2(new_n558_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n493_), .B(new_n502_), .C1(new_n516_), .C2(new_n509_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(new_n208_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n245_), .A2(new_n246_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n562_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT75), .B(new_n562_), .C1(new_n564_), .C2(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n247_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n521_), .A2(new_n232_), .A3(new_n525_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n560_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT72), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n571_), .A2(new_n575_), .A3(new_n572_), .A4(new_n560_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n569_), .A2(new_n570_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n577_), .A2(KEYINPUT73), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n577_), .B2(KEYINPUT73), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT76), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT76), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n569_), .A2(new_n570_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n574_), .A2(new_n576_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT73), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n584_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n577_), .A2(KEYINPUT73), .A3(new_n584_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n582_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT76), .A3(new_n588_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n470_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n244_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n603_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n603_), .A2(new_n609_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n600_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n462_), .A2(new_n555_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT104), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(new_n416_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n456_), .A2(new_n461_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n598_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n614_), .B1(new_n622_), .B2(KEYINPUT105), .ZN(new_n623_));
  INV_X1    g422(.A(new_n555_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n262_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n626_), .A3(new_n598_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n459_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n618_), .A2(new_n619_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n620_), .A2(new_n629_), .A3(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n457_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n617_), .A2(new_n210_), .A3(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n623_), .A2(new_n625_), .A3(new_n632_), .A4(new_n627_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(G8gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n634_), .B2(G8gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n639_), .B(new_n641_), .ZN(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n628_), .B2(new_n315_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT41), .Z(new_n644_));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n617_), .A2(new_n645_), .A3(new_n458_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1326gat));
  OAI21_X1  g446(.A(G22gat), .B1(new_n628_), .B2(new_n460_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n460_), .A2(G22gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT107), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n617_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(G1327gat));
  NAND2_X1  g452(.A1(new_n587_), .A2(new_n614_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n624_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n462_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n416_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n625_), .A2(new_n614_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n621_), .B2(new_n600_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n600_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT43), .B(new_n662_), .C1(new_n456_), .C2(new_n461_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n659_), .B(KEYINPUT44), .C1(new_n661_), .C2(new_n663_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n416_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n657_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT111), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT110), .B1(new_n671_), .B2(KEYINPUT46), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n632_), .A3(new_n667_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n457_), .A2(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n462_), .A2(new_n655_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n462_), .A2(new_n678_), .A3(new_n655_), .A4(new_n675_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(KEYINPUT45), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT45), .B1(new_n677_), .B2(new_n679_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n672_), .B1(new_n674_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n674_), .A2(new_n684_), .A3(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n671_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1329gat));
  NAND3_X1  g487(.A1(new_n668_), .A2(G43gat), .A3(new_n458_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G43gat), .B1(new_n656_), .B2(new_n458_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT112), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n656_), .B2(new_n440_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n440_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n668_), .B2(new_n698_), .ZN(G1331gat));
  INV_X1    g498(.A(new_n262_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n624_), .A3(new_n615_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT113), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OR3_X1    g503(.A1(new_n704_), .A2(G57gat), .A3(new_n459_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n555_), .A2(new_n700_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n623_), .A2(new_n627_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n459_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g508(.A(G64gat), .B1(new_n707_), .B2(new_n457_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n457_), .A2(G64gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n704_), .B2(new_n712_), .ZN(G1333gat));
  OAI21_X1  g512(.A(G71gat), .B1(new_n707_), .B2(new_n315_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n264_), .A3(new_n458_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1334gat));
  OAI21_X1  g516(.A(G78gat), .B1(new_n707_), .B2(new_n460_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT50), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n460_), .A2(G78gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n704_), .B2(new_n720_), .ZN(G1335gat));
  INV_X1    g520(.A(G85gat), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n661_), .A2(new_n663_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n555_), .A2(new_n700_), .A3(new_n613_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n722_), .B1(new_n725_), .B2(new_n416_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n701_), .A2(new_n624_), .A3(new_n587_), .A4(new_n614_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(G85gat), .A3(new_n459_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1336gat));
  NOR3_X1   g528(.A1(new_n727_), .A2(G92gat), .A3(new_n457_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n632_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G92gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1337gat));
  NOR3_X1   g533(.A1(new_n727_), .A2(new_n491_), .A3(new_n315_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n725_), .A2(new_n458_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G99gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1338gat));
  OAI211_X1 g538(.A(new_n440_), .B(new_n724_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n440_), .A2(new_n423_), .ZN(new_n744_));
  OAI22_X1  g543(.A1(new_n742_), .A2(new_n743_), .B1(new_n727_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g545(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n615_), .A2(new_n262_), .A3(new_n555_), .A4(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n555_), .A2(new_n591_), .A3(new_n613_), .A4(new_n599_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n700_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n546_), .A2(new_n550_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n550_), .A2(KEYINPUT56), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n528_), .A2(new_n533_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n544_), .A2(new_n536_), .A3(new_n538_), .A4(new_n518_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n757_), .A2(KEYINPUT55), .B1(new_n758_), .B2(new_n540_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n534_), .A2(new_n760_), .A3(new_n545_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n550_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n755_), .A2(new_n762_), .B1(new_n764_), .B2(KEYINPUT56), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n762_), .A2(new_n755_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n754_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT117), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n754_), .B(new_n769_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n243_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n227_), .B(new_n771_), .C1(new_n244_), .C2(new_n247_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n251_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n252_), .A2(new_n257_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n551_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n768_), .A2(new_n770_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n598_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n546_), .A2(new_n550_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n764_), .A2(KEYINPUT56), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n774_), .B(new_n780_), .C1(new_n781_), .C2(new_n762_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n762_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(KEYINPUT56), .B2(new_n764_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n780_), .A4(new_n774_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n600_), .A2(new_n784_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n591_), .A2(new_n599_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n787_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n587_), .A2(new_n778_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n776_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n779_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n752_), .B1(new_n796_), .B2(new_n614_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n632_), .A2(new_n459_), .A3(new_n440_), .A4(new_n315_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n775_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n767_), .B2(KEYINPUT117), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n587_), .B1(new_n802_), .B2(new_n770_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n795_), .B(new_n788_), .C1(new_n803_), .C2(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n752_), .B1(new_n614_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n800_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n262_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n797_), .A2(new_n799_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n700_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1340gat));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n795_), .B1(new_n803_), .B2(KEYINPUT57), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n791_), .B1(new_n790_), .B2(new_n787_), .ZN(new_n816_));
  AND4_X1   g615(.A1(new_n791_), .A2(new_n600_), .A3(new_n784_), .A4(new_n787_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n614_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n752_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n814_), .B1(new_n821_), .B2(new_n798_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n624_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT120), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n795_), .A2(new_n788_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n776_), .B2(new_n598_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n614_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n820_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n555_), .B1(new_n828_), .B2(new_n806_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n800_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(G120gat), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n555_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n810_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(KEYINPUT121), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n808_), .B2(new_n614_), .ZN(new_n841_));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n810_), .A2(new_n842_), .A3(new_n613_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT122), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1342gat));
  OAI21_X1  g647(.A(G134gat), .B1(new_n808_), .B2(new_n662_), .ZN(new_n849_));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n810_), .A2(new_n850_), .A3(new_n587_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n315_), .A2(new_n440_), .ZN(new_n853_));
  OR4_X1    g652(.A1(new_n459_), .A2(new_n797_), .A3(new_n632_), .A4(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n262_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT123), .B(G141gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n555_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT124), .B(G148gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  NOR2_X1   g659(.A1(new_n854_), .A2(new_n614_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT61), .B(G155gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  OAI21_X1  g662(.A(G162gat), .B1(new_n854_), .B2(new_n662_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n598_), .A2(G162gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n854_), .B2(new_n865_), .ZN(G1347gat));
  NAND4_X1  g665(.A1(new_n632_), .A2(new_n459_), .A3(new_n460_), .A4(new_n458_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n805_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869_), .B2(new_n262_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(KEYINPUT62), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n870_), .A2(KEYINPUT62), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n868_), .A2(new_n700_), .A3(new_n340_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1348gat));
  AOI21_X1  g673(.A(G176gat), .B1(new_n868_), .B2(new_n624_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n797_), .A2(new_n867_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n555_), .A2(new_n290_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  AOI21_X1  g677(.A(G183gat), .B1(new_n876_), .B2(new_n613_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n614_), .A2(new_n282_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n868_), .B2(new_n880_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n869_), .B2(new_n662_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(new_n285_), .A3(new_n587_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1351gat));
  NOR3_X1   g683(.A1(new_n457_), .A2(new_n853_), .A3(new_n416_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n821_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT125), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n700_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT126), .B(G197gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n624_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT127), .B(G204gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1353gat));
  AOI211_X1 g692(.A(KEYINPUT63), .B(G211gat), .C1(new_n887_), .C2(new_n613_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  AND3_X1   g694(.A1(new_n887_), .A2(new_n613_), .A3(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n887_), .A2(new_n898_), .A3(new_n587_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n887_), .A2(new_n600_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1355gat));
endmodule


