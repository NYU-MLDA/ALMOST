//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G15gat), .ZN(new_n206_));
  INV_X1    g005(.A(G15gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G22gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT79), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT79), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G1gat), .B(G8gat), .Z(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n213_), .A3(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G231gat), .A2(G233gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G71gat), .B(G78gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n222_), .B1(KEYINPUT11), .B2(new_n220_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n219_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G155gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT16), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT17), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n230_), .B2(KEYINPUT80), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT34), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT35), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n248_));
  INV_X1    g047(.A(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT65), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n248_), .A2(new_n250_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT9), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G85gat), .A3(G92gat), .ZN(new_n259_));
  INV_X1    g058(.A(G85gat), .ZN(new_n260_));
  INV_X1    g059(.A(G92gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G85gat), .A2(G92gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(KEYINPUT9), .A3(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n254_), .A2(new_n257_), .A3(new_n259_), .A4(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n270_), .A2(new_n259_), .A3(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(KEYINPUT66), .A3(new_n254_), .A4(new_n264_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G99gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n249_), .A3(KEYINPUT67), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT7), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n278_), .A2(new_n275_), .A3(new_n249_), .A4(KEYINPUT67), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n257_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n262_), .A2(new_n263_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(KEYINPUT8), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(KEYINPUT68), .A3(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT8), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n277_), .A2(new_n279_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n270_), .A2(KEYINPUT69), .A3(new_n271_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n281_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n288_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n247_), .B(new_n274_), .C1(new_n287_), .C2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n281_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n285_), .B(new_n286_), .C1(new_n300_), .C2(new_n288_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(KEYINPUT72), .A3(new_n247_), .A4(new_n274_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n274_), .B1(new_n287_), .B2(new_n296_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n247_), .B(KEYINPUT15), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n304_), .A2(new_n305_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n244_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G190gat), .B(G218gat), .Z(new_n309_));
  XOR2_X1   g108(.A(G134gat), .B(G162gat), .Z(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n241_), .A2(new_n242_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n267_), .A2(new_n273_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n280_), .A2(KEYINPUT68), .A3(new_n282_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT68), .B1(new_n280_), .B2(new_n282_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n277_), .A2(new_n279_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT8), .B1(new_n322_), .B2(new_n281_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n245_), .B(new_n246_), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT15), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n316_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n315_), .B1(new_n328_), .B2(new_n244_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n303_), .A2(new_n315_), .A3(new_n244_), .A4(new_n306_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n308_), .B(new_n314_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT37), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n303_), .A2(new_n244_), .A3(new_n306_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT74), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n307_), .B1(new_n335_), .B2(new_n330_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n337_));
  XOR2_X1   g136(.A(new_n311_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n332_), .B(new_n333_), .C1(new_n336_), .C2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT78), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n330_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n308_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT77), .A3(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n332_), .A2(KEYINPUT75), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n336_), .A2(new_n348_), .A3(new_n314_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT37), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n238_), .B1(new_n341_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G230gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT64), .Z(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT70), .B1(new_n304_), .B2(new_n228_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n324_), .A2(new_n356_), .A3(new_n229_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n324_), .A2(new_n229_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n354_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n354_), .B1(new_n324_), .B2(new_n229_), .ZN(new_n361_));
  AOI211_X1 g160(.A(KEYINPUT12), .B(new_n229_), .C1(new_n301_), .C2(new_n274_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT12), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n304_), .B2(new_n228_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n361_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT5), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G176gat), .B(G204gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(new_n365_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT13), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT13), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT71), .B1(new_n375_), .B2(new_n377_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G155gat), .ZN(new_n384_));
  INV_X1    g183(.A(G162gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT89), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(G155gat), .B2(G162gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n390_), .A2(KEYINPUT1), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n389_), .A2(new_n390_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT102), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n396_), .A2(new_n400_), .B1(new_n402_), .B2(new_n409_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT102), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G127gat), .B(G134gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n413_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT0), .ZN(new_n426_));
  INV_X1    g225(.A(G57gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G85gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n411_), .A2(new_n430_), .A3(new_n418_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n423_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n424_), .B(new_n429_), .C1(new_n431_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT103), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n429_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n424_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n431_), .A2(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n436_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G211gat), .B(G218gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445_));
  INV_X1    g244(.A(G197gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(G204gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(KEYINPUT21), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G197gat), .B(G204gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(KEYINPUT21), .A3(new_n444_), .A4(new_n447_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n444_), .A2(KEYINPUT21), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT24), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT100), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT86), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n464_), .A3(KEYINPUT23), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G183gat), .A3(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(KEYINPUT25), .B(G183gat), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT26), .B(G190gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n460_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT22), .B(G169gat), .Z(new_n475_));
  OAI21_X1  g274(.A(new_n456_), .B1(new_n475_), .B2(G176gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n461_), .A2(KEYINPUT23), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT85), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n462_), .A2(new_n464_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT87), .B1(new_n479_), .B2(new_n466_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n481_), .B(KEYINPUT23), .C1(new_n462_), .C2(new_n464_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n478_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G183gat), .A2(G190gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n455_), .B1(new_n474_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n484_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n476_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n489_), .B2(new_n488_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(KEYINPUT82), .A3(G183gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n470_), .B2(KEYINPUT82), .ZN(new_n494_));
  INV_X1    g293(.A(G190gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT83), .B1(new_n495_), .B2(KEYINPUT26), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n494_), .B(new_n496_), .C1(KEYINPUT83), .C2(new_n472_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n457_), .A2(KEYINPUT84), .A3(new_n459_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT84), .B1(new_n457_), .B2(new_n459_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n469_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n483_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n501_), .A3(new_n454_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n487_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n503_), .A2(KEYINPUT20), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n491_), .A2(new_n501_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n508_), .B2(new_n454_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT99), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT99), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(KEYINPUT20), .C1(new_n508_), .C2(new_n454_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n454_), .B1(new_n474_), .B2(new_n486_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n506_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n507_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G8gat), .B(G36gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT18), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G64gat), .B(G92gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT32), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n503_), .A2(KEYINPUT20), .A3(new_n515_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n514_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n515_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n443_), .B(new_n522_), .C1(new_n525_), .C2(new_n521_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n520_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n514_), .A2(new_n515_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT101), .B(new_n527_), .C1(new_n528_), .C2(new_n507_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT101), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n516_), .A2(new_n520_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n435_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n435_), .A2(new_n534_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n429_), .B1(new_n433_), .B2(new_n422_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n432_), .A2(new_n423_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n431_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n526_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G22gat), .B(G50gat), .Z(new_n542_));
  NOR3_X1   g341(.A1(new_n411_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n413_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n542_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT28), .B1(new_n411_), .B2(KEYINPUT29), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n413_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n542_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT91), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT94), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n454_), .B1(new_n413_), .B2(new_n545_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(KEYINPUT92), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n454_), .B(KEYINPUT94), .C1(new_n413_), .C2(new_n545_), .ZN(new_n559_));
  INV_X1    g358(.A(G228gat), .ZN(new_n560_));
  INV_X1    g359(.A(G233gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  OAI221_X1 g362(.A(new_n556_), .B1(new_n560_), .B2(new_n561_), .C1(new_n557_), .C2(KEYINPUT92), .ZN(new_n564_));
  XOR2_X1   g363(.A(G78gat), .B(G106gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT95), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT96), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n563_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n553_), .B(new_n555_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n564_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n573_), .A2(new_n551_), .A3(new_n547_), .A4(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n570_), .A2(new_n575_), .A3(KEYINPUT97), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G71gat), .B(G99gat), .ZN(new_n577_));
  INV_X1    g376(.A(G43gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G227gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n207_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n579_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n491_), .A2(new_n501_), .A3(KEYINPUT30), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT30), .B1(new_n491_), .B2(new_n501_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n418_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT31), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n419_), .A3(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT97), .B1(new_n570_), .B2(new_n575_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n576_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n541_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n443_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n593_), .A2(new_n597_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n576_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n553_), .A2(new_n555_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n563_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n573_), .B2(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n609_), .A2(new_n569_), .A3(new_n552_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n570_), .A2(new_n575_), .A3(KEYINPUT97), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n611_), .A2(new_n612_), .B1(new_n597_), .B2(new_n593_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n602_), .B1(new_n604_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT27), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n533_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n516_), .A2(new_n520_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n527_), .B(new_n523_), .C1(new_n524_), .C2(new_n515_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT27), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n601_), .B1(new_n614_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n217_), .A2(new_n305_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n215_), .A2(new_n216_), .A3(new_n247_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n216_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n213_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n325_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n625_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n623_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT81), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n626_), .A2(new_n631_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n634_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n631_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n630_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n636_), .B(new_n638_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n635_), .B1(new_n639_), .B2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n352_), .A2(new_n383_), .A3(new_n621_), .A4(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT104), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n602_), .A2(G1gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n603_), .B1(new_n576_), .B2(new_n599_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n598_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n443_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n619_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n533_), .B2(new_n615_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n652_), .A2(new_n654_), .B1(new_n541_), .B2(new_n600_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n644_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n378_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n339_), .B1(new_n342_), .B2(new_n308_), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n307_), .B(new_n313_), .C1(new_n335_), .C2(new_n330_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT105), .Z(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n238_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n602_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n649_), .A2(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n658_), .A2(new_n663_), .A3(new_n620_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n669_), .B2(KEYINPUT39), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n668_), .A2(KEYINPUT106), .A3(new_n671_), .A4(G8gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(KEYINPUT39), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n646_), .A2(new_n203_), .A3(new_n620_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n675_), .A3(KEYINPUT40), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n664_), .B2(new_n603_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n683_));
  INV_X1    g482(.A(new_n645_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n207_), .A3(new_n598_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n576_), .A2(new_n599_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G22gat), .B1(new_n664_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n687_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n684_), .A2(new_n205_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1327gat));
  INV_X1    g492(.A(new_n661_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n237_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n658_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n443_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n657_), .A2(new_n237_), .A3(new_n656_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT78), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n340_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n661_), .A2(KEYINPUT78), .A3(new_n333_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n351_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n655_), .A2(new_n702_), .A3(KEYINPUT43), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n350_), .A2(KEYINPUT37), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n700_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n621_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n698_), .B1(new_n703_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(G29gat), .A3(new_n443_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT44), .B(new_n698_), .C1(new_n703_), .C2(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  INV_X1    g513(.A(new_n698_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n655_), .B2(new_n702_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n621_), .A2(new_n707_), .A3(new_n704_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n697_), .B1(new_n712_), .B2(new_n721_), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n620_), .B1(new_n718_), .B2(KEYINPUT44), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n721_), .B2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n658_), .A2(new_n724_), .A3(new_n620_), .A4(new_n695_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT45), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n723_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n725_), .B1(new_n714_), .B2(new_n720_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT46), .B(new_n729_), .C1(new_n732_), .C2(new_n724_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1329gat));
  XOR2_X1   g533(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n735_));
  NOR2_X1   g534(.A1(new_n603_), .A2(new_n578_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n711_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n714_), .B2(new_n720_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G43gat), .B1(new_n696_), .B2(new_n598_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n721_), .A2(new_n711_), .A3(new_n736_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n739_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n735_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n740_), .A2(new_n744_), .ZN(G1330gat));
  NOR2_X1   g544(.A1(new_n687_), .A2(G50gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT111), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n696_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n687_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n721_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n721_), .B2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n657_), .A2(KEYINPUT71), .ZN(new_n755_));
  INV_X1    g554(.A(new_n381_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n656_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n655_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n663_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n427_), .A3(new_n602_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n378_), .A2(new_n644_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n352_), .A2(new_n621_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n602_), .B1(new_n762_), .B2(KEYINPUT112), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(KEYINPUT112), .B2(new_n762_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n764_), .B2(new_n427_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT113), .Z(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n759_), .B2(new_n654_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n654_), .A2(G64gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n762_), .B2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n759_), .B2(new_n603_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n603_), .A2(G71gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n762_), .B2(new_n773_), .ZN(G1334gat));
  OAI21_X1  g573(.A(G78gat), .B1(new_n759_), .B2(new_n687_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n687_), .A2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n762_), .B2(new_n777_), .ZN(G1335gat));
  NAND3_X1  g577(.A1(new_n758_), .A2(KEYINPUT114), .A3(new_n695_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n380_), .A2(new_n381_), .A3(new_n644_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n621_), .A2(new_n695_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n260_), .B1(new_n785_), .B2(new_n602_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n761_), .A2(new_n238_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n443_), .A2(G85gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT116), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n787_), .A2(new_n788_), .B1(new_n790_), .B2(new_n792_), .ZN(G1336gat));
  AOI21_X1  g592(.A(G92gat), .B1(new_n784_), .B2(new_n620_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n620_), .A2(G92gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT117), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n790_), .B2(new_n796_), .ZN(G1337gat));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n598_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n598_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n799_), .A2(G99gat), .B1(new_n784_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT114), .B1(new_n758_), .B2(new_n695_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n781_), .A2(new_n782_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n603_), .B(new_n789_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n806_), .B(new_n798_), .C1(new_n807_), .C2(new_n275_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT51), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n803_), .A2(new_n809_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n798_), .B(KEYINPUT51), .C1(new_n801_), .C2(new_n802_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1338gat));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n790_), .A2(new_n691_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G106gat), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT52), .B(new_n249_), .C1(new_n790_), .C2(new_n691_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n691_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n815_), .A2(new_n816_), .B1(new_n785_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  OAI221_X1 g619(.A(new_n820_), .B1(new_n785_), .B2(new_n817_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  NAND2_X1  g621(.A1(new_n654_), .A2(new_n443_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n604_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n644_), .A2(new_n373_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n362_), .A2(new_n364_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n354_), .B1(new_n827_), .B2(new_n358_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n365_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT55), .B(new_n361_), .C1(new_n362_), .C2(new_n364_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n370_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n370_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n826_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT81), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n642_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n630_), .B1(new_n629_), .B2(new_n623_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n638_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n638_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n844_), .B(new_n845_), .C1(new_n625_), .C2(new_n624_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n374_), .A2(new_n840_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n694_), .B1(new_n837_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n366_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n851_), .A2(new_n372_), .B1(new_n840_), .B2(new_n635_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n370_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n370_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n374_), .A2(new_n840_), .A3(new_n846_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT57), .A3(new_n694_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n840_), .A2(new_n373_), .A3(new_n846_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT121), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(KEYINPUT121), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n859_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n850_), .B(new_n858_), .C1(new_n702_), .C2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n657_), .A2(new_n644_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(new_n237_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n866_), .A2(new_n238_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n867_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n825_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n644_), .ZN(new_n875_));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n825_), .C1(new_n870_), .C2(new_n872_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n857_), .B2(new_n694_), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n849_), .B(new_n661_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n341_), .A2(new_n351_), .A3(new_n862_), .A4(new_n864_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n237_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT54), .B1(new_n352_), .B2(new_n868_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n884_), .A2(new_n871_), .A3(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n879_), .B(KEYINPUT59), .C1(new_n886_), .C2(new_n825_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n656_), .B(new_n876_), .C1(new_n878_), .C2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n875_), .B1(new_n888_), .B2(new_n874_), .ZN(G1340gat));
  NOR3_X1   g688(.A1(new_n378_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n873_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n383_), .B(new_n876_), .C1(new_n878_), .C2(new_n887_), .ZN(new_n893_));
  INV_X1    g692(.A(G120gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1341gat));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n873_), .A2(new_n896_), .A3(new_n237_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n238_), .B(new_n876_), .C1(new_n878_), .C2(new_n887_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1342gat));
  XNOR2_X1  g698(.A(KEYINPUT124), .B(G134gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n707_), .A2(new_n900_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n901_), .B(new_n876_), .C1(new_n878_), .C2(new_n887_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n662_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n886_), .A2(new_n903_), .A3(new_n825_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n904_), .B2(G134gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n873_), .A2(new_n662_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  INV_X1    g706(.A(G134gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n902_), .A2(new_n910_), .ZN(G1343gat));
  NOR2_X1   g710(.A1(new_n886_), .A2(new_n650_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(new_n644_), .A3(new_n824_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n382_), .A3(new_n824_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n237_), .A3(new_n824_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  NOR2_X1   g718(.A1(new_n903_), .A2(G162gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n824_), .A3(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n870_), .A2(new_n872_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n922_), .A2(new_n613_), .A3(new_n707_), .A4(new_n824_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G162gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n921_), .A2(new_n924_), .A3(KEYINPUT125), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n654_), .A2(new_n443_), .A3(new_n651_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n922_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n644_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n933_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n931_), .A2(new_n656_), .ZN(new_n936_));
  INV_X1    g735(.A(G169gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n934_), .B(new_n938_), .C1(new_n475_), .C2(new_n933_), .ZN(G1348gat));
  OR3_X1    g738(.A1(new_n931_), .A2(G176gat), .A3(new_n378_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G176gat), .B1(new_n931_), .B2(new_n383_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n931_), .A2(new_n238_), .ZN(new_n943_));
  MUX2_X1   g742(.A(G183gat), .B(new_n471_), .S(new_n943_), .Z(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n931_), .B2(new_n702_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n662_), .A2(new_n472_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n931_), .B2(new_n946_), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n654_), .A2(new_n443_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n912_), .A2(new_n644_), .A3(new_n948_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g749(.A1(new_n912_), .A2(new_n382_), .A3(new_n948_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g751(.A1(new_n922_), .A2(new_n237_), .A3(new_n613_), .A4(new_n948_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955_));
  INV_X1    g754(.A(G211gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT126), .B1(new_n954_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n953_), .A2(new_n959_), .A3(new_n955_), .A4(new_n956_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT63), .B(G211gat), .Z(new_n961_));
  AOI22_X1  g760(.A1(new_n958_), .A2(new_n960_), .B1(new_n954_), .B2(new_n961_), .ZN(G1354gat));
  AND4_X1   g761(.A1(new_n662_), .A2(new_n922_), .A3(new_n613_), .A4(new_n948_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964_));
  OR2_X1    g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(G218gat), .B1(new_n963_), .B2(new_n964_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n912_), .A2(new_n948_), .ZN(new_n967_));
  AND2_X1   g766(.A1(new_n707_), .A2(G218gat), .ZN(new_n968_));
  AOI22_X1  g767(.A1(new_n965_), .A2(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(G1355gat));
endmodule


