//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_;
  XOR2_X1   g000(.A(KEYINPUT26), .B(G190gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203_));
  INV_X1    g002(.A(G183gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT25), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT88), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G183gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n203_), .B(new_n206_), .C1(new_n209_), .C2(KEYINPUT88), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n208_), .A2(KEYINPUT88), .A3(new_n203_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n202_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n214_), .B(new_n219_), .C1(KEYINPUT24), .C2(new_n217_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n218_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n216_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n223_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G113gat), .ZN(new_n233_));
  INV_X1    g032(.A(G120gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT31), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n244_), .A3(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT95), .ZN(new_n254_));
  INV_X1    g053(.A(G204gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G197gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT94), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT96), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n251_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n260_), .B(KEYINPUT21), .C1(new_n259_), .C2(new_n258_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n256_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT21), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n251_), .B(new_n263_), .C1(new_n258_), .C2(KEYINPUT21), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n266_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268_));
  OAI221_X1 g067(.A(new_n267_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(KEYINPUT92), .Z(new_n270_));
  NOR2_X1   g069(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n271_));
  INV_X1    g070(.A(G141gat), .ZN(new_n272_));
  INV_X1    g071(.A(G148gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NOR4_X1   g073(.A1(KEYINPUT91), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT2), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n276_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n278_));
  NOR4_X1   g077(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n269_), .B1(new_n270_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT29), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n265_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G78gat), .B(G106gat), .Z(new_n285_));
  AOI21_X1  g084(.A(new_n250_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n284_), .A2(KEYINPUT97), .A3(new_n285_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT93), .A3(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n280_), .A2(KEYINPUT29), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G22gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT28), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT93), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n287_), .A2(new_n295_), .A3(new_n288_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT98), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n284_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n284_), .A2(new_n298_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n293_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n235_), .B(new_n280_), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT4), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n235_), .A2(new_n308_), .A3(new_n280_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT103), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT103), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n304_), .A2(new_n306_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G57gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G85gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT104), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT33), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(KEYINPUT33), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n304_), .A2(new_n307_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n305_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n317_), .B(new_n323_), .C1(new_n324_), .C2(new_n307_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n261_), .A2(new_n264_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n202_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n220_), .B1(new_n328_), .B2(new_n209_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n227_), .B2(new_n222_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT99), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT19), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  INV_X1    g134(.A(new_n230_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n327_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n327_), .A2(new_n330_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n339_), .B(KEYINPUT20), .C1(new_n336_), .C2(new_n327_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G8gat), .B(G36gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT101), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  OR3_X1    g148(.A1(new_n343_), .A2(KEYINPUT102), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n349_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n352_), .A3(new_n342_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(KEYINPUT102), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n326_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n332_), .A2(new_n341_), .A3(new_n337_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n340_), .A2(new_n334_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n312_), .A2(new_n313_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n317_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n361_), .A2(new_n319_), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n359_), .B(new_n362_), .C1(new_n343_), .C2(new_n356_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n249_), .B(new_n303_), .C1(new_n355_), .C2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n303_), .A2(new_n248_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n294_), .A2(new_n302_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n354_), .A2(new_n350_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT107), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT107), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n354_), .A2(new_n350_), .A3(new_n371_), .A4(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT106), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n351_), .B(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n352_), .A2(KEYINPUT105), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n352_), .A2(KEYINPUT105), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n368_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n367_), .A2(new_n370_), .A3(new_n372_), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n362_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n364_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G29gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G43gat), .B(G50gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n383_), .B(new_n384_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n386_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G22gat), .ZN(new_n392_));
  INV_X1    g191(.A(G1gat), .ZN(new_n393_));
  INV_X1    g192(.A(G8gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT14), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G8gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n391_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT84), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G229gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT85), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n391_), .B(KEYINPUT15), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n401_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n400_), .A2(new_n409_), .A3(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G113gat), .B(G141gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(new_n215_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(new_n252_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .A4(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n417_), .A2(KEYINPUT86), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(KEYINPUT86), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n415_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n417_), .B(KEYINPUT86), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(KEYINPUT87), .A3(new_n415_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G57gat), .B(G64gat), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n428_), .A2(KEYINPUT11), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(KEYINPUT11), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G71gat), .B(G78gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT73), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n440_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  NOR2_X1   g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT67), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT7), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT68), .B1(new_n456_), .B2(new_n449_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n446_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n439_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n448_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(KEYINPUT68), .A3(new_n449_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n445_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n468_), .A2(KEYINPUT69), .A3(new_n463_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n441_), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT70), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT71), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n440_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n472_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n477_), .B(new_n481_), .C1(new_n451_), .C2(new_n457_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n462_), .B1(new_n482_), .B2(new_n461_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n438_), .B1(new_n470_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n458_), .A2(new_n439_), .A3(new_n464_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT69), .B1(new_n468_), .B2(new_n463_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n461_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n489_), .A3(KEYINPUT72), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT64), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT65), .B(G106gat), .Z(new_n494_));
  OAI21_X1  g293(.A(new_n479_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n460_), .A2(KEYINPUT66), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n496_), .B(KEYINPUT9), .Z(new_n497_));
  AND2_X1   g296(.A1(new_n497_), .A2(new_n459_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n437_), .B1(new_n491_), .B2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n487_), .A2(new_n489_), .A3(KEYINPUT72), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT72), .B1(new_n487_), .B2(new_n489_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n437_), .B(new_n500_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n436_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n434_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G230gat), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n507_), .B2(new_n434_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n434_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n511_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G120gat), .B(G148gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G176gat), .B(G204gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT76), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n514_), .A2(new_n526_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n523_), .B(KEYINPUT75), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT77), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT77), .ZN(new_n534_));
  AOI211_X1 g333(.A(new_n534_), .B(new_n531_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT13), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT73), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n504_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n509_), .B1(new_n539_), .B2(new_n436_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n517_), .B1(new_n540_), .B2(new_n513_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n526_), .B1(new_n541_), .B2(new_n523_), .ZN(new_n542_));
  AND4_X1   g341(.A1(new_n526_), .A2(new_n514_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n532_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n534_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n528_), .A2(KEYINPUT77), .A3(new_n532_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n426_), .B1(new_n536_), .B2(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n382_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n539_), .A2(new_n406_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n507_), .A2(new_n391_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(KEYINPUT35), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n552_), .A2(new_n559_), .A3(new_n560_), .A4(new_n553_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G134gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(G162gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n561_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT36), .A3(new_n565_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT81), .ZN(new_n572_));
  OR3_X1    g371(.A1(new_n571_), .A2(new_n572_), .A3(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n398_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n434_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT82), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT16), .B(G183gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT83), .Z(new_n590_));
  INV_X1    g389(.A(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n587_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n578_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n551_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n393_), .A3(new_n381_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n571_), .A2(new_n594_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n550_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n362_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n370_), .A2(new_n372_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n379_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n550_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G8gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n611_), .A3(G8gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT109), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n597_), .A2(new_n394_), .A3(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n605_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT40), .A3(new_n616_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n602_), .B2(new_n249_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(G15gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n597_), .A2(new_n626_), .A3(new_n248_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT110), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1326gat));
  OAI21_X1  g429(.A(G22gat), .B1(new_n602_), .B2(new_n303_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  INV_X1    g431(.A(G22gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n303_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n597_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1327gat));
  NAND2_X1  g435(.A1(new_n571_), .A2(new_n594_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT112), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n550_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n381_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n577_), .A2(new_n382_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT111), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n577_), .A2(new_n382_), .A3(new_n645_), .A4(KEYINPUT43), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n594_), .A3(new_n549_), .A4(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n362_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n642_), .B1(new_n653_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n641_), .A2(new_n655_), .A3(new_n607_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT45), .ZN(new_n657_));
  INV_X1    g456(.A(new_n607_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n651_), .A2(new_n652_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(new_n655_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n657_), .B(KEYINPUT46), .C1(new_n659_), .C2(new_n655_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  XOR2_X1   g463(.A(KEYINPUT113), .B(G43gat), .Z(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n641_), .B2(new_n248_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n649_), .B(KEYINPUT44), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n248_), .A2(G43gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1330gat));
  AOI21_X1  g470(.A(G50gat), .B1(new_n641_), .B2(new_n634_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n634_), .A2(G50gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n667_), .B2(new_n673_), .ZN(G1331gat));
  NAND2_X1  g473(.A1(new_n536_), .A2(new_n548_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n425_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n382_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(new_n594_), .A3(new_n571_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(G57gat), .A3(new_n381_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT114), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT114), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n596_), .A2(new_n677_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n362_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n680_), .B(new_n681_), .C1(G57gat), .C2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT115), .Z(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n678_), .B2(new_n607_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT48), .Z(new_n688_));
  INV_X1    g487(.A(new_n682_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n686_), .A3(new_n607_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1333gat));
  INV_X1    g490(.A(G71gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n678_), .B2(new_n248_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT49), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n692_), .A3(new_n248_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n678_), .B2(new_n634_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT50), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n697_), .A3(new_n634_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1335gat));
  NAND3_X1  g500(.A1(new_n639_), .A2(new_n382_), .A3(new_n676_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n381_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n647_), .A2(new_n594_), .A3(new_n648_), .A4(new_n676_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n362_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n706_), .B2(G85gat), .ZN(G1336gat));
  NAND2_X1  g506(.A1(new_n607_), .A2(G92gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT116), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n702_), .A2(new_n658_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n705_), .A2(new_n709_), .B1(new_n710_), .B2(G92gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT117), .ZN(G1337gat));
  OAI21_X1  g511(.A(G99gat), .B1(new_n705_), .B2(new_n249_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n249_), .A2(new_n493_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n702_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g515(.A(G106gat), .B1(new_n705_), .B2(new_n303_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT52), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n719_), .B(G106gat), .C1(new_n705_), .C2(new_n303_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n702_), .A2(new_n494_), .A3(new_n303_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT53), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  NOR2_X1   g526(.A1(new_n607_), .A2(new_n362_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n248_), .A3(new_n303_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT122), .Z(new_n730_));
  INV_X1    g529(.A(new_n571_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n506_), .A2(new_n516_), .A3(new_n510_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n512_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n514_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n540_), .A2(KEYINPUT55), .A3(new_n513_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n529_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT120), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT120), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n741_), .A3(new_n529_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT121), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n529_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n739_), .A2(KEYINPUT121), .A3(new_n740_), .A4(new_n742_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n425_), .A2(new_n528_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n545_), .A2(new_n547_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n400_), .A2(new_n401_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n407_), .A2(new_n402_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n414_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n423_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT57), .B(new_n731_), .C1(new_n750_), .C2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n748_), .A2(new_n749_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n571_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n738_), .A2(new_n740_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n746_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n528_), .A3(new_n755_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT58), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n577_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(new_n760_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n594_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n675_), .A2(new_n595_), .A3(new_n426_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n425_), .B1(new_n536_), .B2(new_n548_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT118), .A3(new_n595_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n769_), .B1(new_n775_), .B2(new_n578_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n577_), .B(new_n768_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n730_), .B1(new_n767_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779_), .B2(new_n425_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  AND4_X1   g580(.A1(KEYINPUT118), .A2(new_n675_), .A3(new_n595_), .A4(new_n426_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT118), .B1(new_n773_), .B2(new_n595_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n578_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n768_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n775_), .A2(new_n578_), .A3(new_n769_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n594_), .B2(new_n766_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n781_), .B1(new_n788_), .B2(new_n730_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n779_), .A2(KEYINPUT59), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n426_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n780_), .B1(new_n791_), .B2(G113gat), .ZN(G1340gat));
  NAND2_X1  g591(.A1(new_n767_), .A2(new_n778_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n730_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n234_), .A2(KEYINPUT60), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n234_), .B1(new_n675_), .B2(KEYINPUT60), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT123), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT124), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT124), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n779_), .A2(new_n800_), .A3(new_n795_), .A4(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n675_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n234_), .ZN(G1341gat));
  AOI21_X1  g603(.A(G127gat), .B1(new_n779_), .B2(new_n595_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n594_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g606(.A(G134gat), .B1(new_n779_), .B2(new_n571_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n578_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n788_), .A2(new_n366_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n425_), .A3(new_n728_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G141gat), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n811_), .A2(new_n272_), .A3(new_n425_), .A4(new_n728_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1344gat));
  INV_X1    g614(.A(new_n675_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n816_), .A3(new_n728_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G148gat), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n811_), .A2(new_n273_), .A3(new_n816_), .A4(new_n728_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1345gat));
  INV_X1    g619(.A(new_n366_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n793_), .A2(new_n595_), .A3(new_n821_), .A4(new_n728_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1346gat));
  NAND4_X1  g623(.A1(new_n811_), .A2(G162gat), .A3(new_n577_), .A4(new_n728_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n793_), .A2(new_n571_), .A3(new_n821_), .A4(new_n728_), .ZN(new_n826_));
  INV_X1    g625(.A(G162gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1347gat));
  NOR3_X1   g628(.A1(new_n658_), .A2(new_n381_), .A3(new_n365_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n793_), .A2(new_n425_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n215_), .B1(new_n832_), .B2(KEYINPUT62), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(KEYINPUT62), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n831_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n793_), .A2(new_n830_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n425_), .A2(new_n226_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT126), .Z(new_n839_));
  OAI22_X1  g638(.A1(new_n835_), .A2(new_n836_), .B1(new_n837_), .B2(new_n839_), .ZN(G1348gat));
  NOR2_X1   g639(.A1(new_n837_), .A2(new_n675_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n216_), .ZN(G1349gat));
  NAND3_X1  g641(.A1(new_n793_), .A2(new_n595_), .A3(new_n830_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n209_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n204_), .B2(new_n843_), .ZN(G1350gat));
  OAI21_X1  g644(.A(G190gat), .B1(new_n837_), .B2(new_n578_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n571_), .A2(new_n328_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n837_), .B2(new_n847_), .ZN(G1351gat));
  NOR2_X1   g647(.A1(new_n658_), .A2(new_n381_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n821_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n767_), .B2(new_n778_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n425_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n816_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g654(.A(KEYINPUT63), .B(G211gat), .C1(new_n851_), .C2(new_n595_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n788_), .A2(new_n594_), .A3(new_n850_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT63), .B(G211gat), .Z(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1354gat));
  AND2_X1   g658(.A1(new_n577_), .A2(G218gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n851_), .A2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n788_), .A2(new_n731_), .A3(new_n850_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT127), .B(new_n861_), .C1(new_n862_), .C2(G218gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT127), .ZN(new_n864_));
  AOI21_X1  g663(.A(G218gat), .B1(new_n851_), .B2(new_n571_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n850_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n793_), .A2(new_n866_), .A3(new_n860_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n868_), .ZN(G1355gat));
endmodule


