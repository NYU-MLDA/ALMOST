//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  INV_X1    g003(.A(G43gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G29gat), .ZN(new_n208_));
  INV_X1    g007(.A(G29gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G36gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n210_), .A3(new_n205_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n206_), .A2(new_n211_), .A3(KEYINPUT71), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G43gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n204_), .A2(new_n205_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G50gat), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n212_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT71), .B1(new_n206_), .B2(new_n211_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n216_), .A3(new_n213_), .ZN(new_n221_));
  AOI21_X1  g020(.A(G50gat), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n203_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n218_), .B1(new_n212_), .B2(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(G50gat), .A3(new_n221_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT15), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G85gat), .B(G92gat), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n229_), .A2(new_n232_), .A3(new_n234_), .A4(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n241_));
  OR3_X1    g040(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT65), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n241_), .B1(new_n247_), .B2(new_n228_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n242_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n246_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n228_), .B(new_n241_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n240_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT68), .ZN(new_n254_));
  INV_X1    g053(.A(new_n240_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n228_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n257_), .B2(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n227_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n258_), .A2(KEYINPUT72), .A3(new_n225_), .A4(new_n224_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n224_), .A2(new_n225_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n253_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT34), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT73), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT36), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n262_), .A2(new_n265_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n273_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n261_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n279_), .B(KEYINPUT36), .Z(new_n287_));
  INV_X1    g086(.A(new_n283_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n281_), .B2(new_n261_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(new_n287_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n202_), .B1(new_n286_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n284_), .B(KEYINPUT74), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT37), .A3(new_n290_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G155gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT16), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G22gat), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  XOR2_X1   g113(.A(G71gat), .B(G78gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G64gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n315_), .B1(KEYINPUT11), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT67), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(KEYINPUT11), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n315_), .B(new_n320_), .C1(KEYINPUT11), .C2(new_n316_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n314_), .B(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n305_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n303_), .B(KEYINPUT17), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n325_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n298_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT76), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G169gat), .ZN(new_n344_));
  INV_X1    g143(.A(G176gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n334_), .A2(new_n338_), .A3(KEYINPUT82), .A4(new_n335_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n350_), .A2(G169gat), .A3(G176gat), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT81), .B1(new_n352_), .B2(new_n345_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n349_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n345_), .A3(KEYINPUT81), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n350_), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT24), .A4(new_n342_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n334_), .A2(new_n335_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n354_), .A2(new_n357_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n348_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT30), .ZN(new_n364_));
  AND2_X1   g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT31), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT83), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT84), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n377_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n373_), .B(new_n379_), .C1(KEYINPUT84), .C2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G197gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G204gat), .ZN(new_n385_));
  INV_X1    g184(.A(G204gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G197gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT21), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n386_), .B2(G197gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n384_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n387_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(KEYINPUT21), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n390_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n388_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n396_), .A2(KEYINPUT90), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n404_), .B2(new_n399_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT87), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT87), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  AND2_X1   g212(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n421_), .A2(G155gat), .A3(G162gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(G155gat), .B2(G162gat), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n423_), .A2(new_n424_), .B1(G155gat), .B2(G162gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n428_), .B(new_n429_), .C1(new_n430_), .C2(new_n422_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G141gat), .B(G148gat), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n407_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G228gat), .ZN(new_n435_));
  INV_X1    g234(.A(G233gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n406_), .A2(new_n438_), .A3(KEYINPUT91), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n396_), .B2(new_n400_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n404_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n420_), .A2(new_n425_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n444_), .A2(new_n407_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n440_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n396_), .A2(new_n400_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n437_), .B1(new_n434_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n437_), .C1(new_n434_), .C2(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT93), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n407_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT88), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(KEYINPUT88), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G22gat), .B(G50gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT28), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n461_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n447_), .A2(new_n453_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n454_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n456_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n464_), .A3(new_n470_), .A4(new_n456_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G57gat), .B(G85gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n426_), .A2(new_n433_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n376_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(KEYINPUT4), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n426_), .A2(new_n376_), .A3(new_n433_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n376_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n486_), .B1(new_n489_), .B2(KEYINPUT4), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n444_), .A2(new_n376_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n483_), .A2(new_n486_), .A3(new_n491_), .A4(KEYINPUT4), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n480_), .B(new_n485_), .C1(new_n490_), .C2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n483_), .A2(new_n479_), .A3(new_n491_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT98), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n478_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G64gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n502_), .A2(G64gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n499_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n502_), .A2(G64gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G92gat), .A3(new_n503_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n441_), .A2(new_n363_), .A3(new_n442_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n337_), .A2(KEYINPUT26), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G190gat), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT94), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT94), .B1(new_n511_), .B2(new_n513_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT25), .B(G183gat), .Z(new_n516_));
  NOR3_X1   g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n354_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT95), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n339_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n334_), .A2(new_n338_), .A3(KEYINPUT95), .A4(new_n335_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n346_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n448_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND4_X1   g326(.A1(KEYINPUT20), .A2(new_n510_), .A3(new_n524_), .A4(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n363_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n404_), .A2(new_n399_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n527_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n509_), .B1(new_n528_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT20), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n363_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n526_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n510_), .A2(new_n524_), .A3(KEYINPUT20), .A4(new_n527_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n540_), .A2(new_n508_), .A3(new_n506_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT27), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n494_), .A2(new_n478_), .A3(new_n496_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n527_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n510_), .A2(new_n524_), .A3(KEYINPUT20), .A4(new_n526_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n509_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n549_), .A3(KEYINPUT27), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n498_), .A2(new_n545_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n383_), .A2(new_n472_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553_));
  AND4_X1   g352(.A1(new_n470_), .A2(new_n467_), .A3(new_n456_), .A4(new_n464_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n457_), .A2(new_n464_), .B1(new_n467_), .B2(new_n456_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n489_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n477_), .B1(new_n558_), .B2(new_n479_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n483_), .A2(KEYINPUT4), .A3(new_n491_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT96), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n484_), .B1(new_n561_), .B2(new_n492_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n562_), .B2(new_n479_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n543_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n546_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n494_), .A2(KEYINPUT33), .A3(new_n478_), .A4(new_n496_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n506_), .A2(KEYINPUT32), .A3(new_n508_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n528_), .A2(new_n535_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n547_), .A2(new_n569_), .A3(new_n548_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n547_), .A2(new_n569_), .A3(KEYINPUT99), .A4(new_n548_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n546_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n497_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n556_), .ZN(new_n579_));
  AND4_X1   g378(.A1(new_n498_), .A2(new_n545_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT100), .A3(new_n472_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n557_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n552_), .B1(new_n582_), .B2(new_n383_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT12), .B1(new_n324_), .B2(new_n253_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n324_), .A2(new_n253_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n260_), .A2(new_n254_), .A3(KEYINPUT12), .A4(new_n324_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n585_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n324_), .A2(new_n253_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n386_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT5), .B(G176gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n593_), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT13), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT69), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G113gat), .B(G141gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT79), .B(G197gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT78), .B(G169gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n264_), .A2(new_n312_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n312_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n224_), .A2(new_n617_), .A3(new_n225_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n227_), .A2(new_n312_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n615_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT77), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n614_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n617_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n621_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT77), .B1(new_n627_), .B2(new_n619_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n615_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n618_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n617_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(new_n614_), .C1(new_n626_), .C2(new_n621_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT80), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n620_), .A2(new_n622_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n632_), .A4(new_n614_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n625_), .A2(new_n628_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n583_), .A2(new_n609_), .A3(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n331_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n576_), .A2(new_n497_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n307_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n296_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n329_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n639_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n641_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n643_), .A2(new_n644_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n545_), .A2(new_n550_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n640_), .A2(new_n308_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G8gat), .B1(new_n649_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(KEYINPUT101), .A2(KEYINPUT39), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n654_), .B(new_n658_), .C1(new_n656_), .C2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(G1325gat));
  NAND2_X1  g461(.A1(new_n331_), .A2(new_n639_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n663_), .A2(G15gat), .A3(new_n383_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT102), .Z(new_n665_));
  OAI21_X1  g464(.A(G15gat), .B1(new_n649_), .B2(new_n383_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT41), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n649_), .B2(new_n556_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n556_), .A2(G22gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n663_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n646_), .A2(new_n328_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT103), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n639_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n642_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n609_), .A2(new_n638_), .A3(new_n328_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n582_), .A2(new_n383_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n552_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n681_), .B2(new_n298_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n295_), .A2(new_n297_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n583_), .A2(new_n683_), .A3(KEYINPUT43), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n677_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n677_), .C1(new_n682_), .C2(new_n684_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n641_), .A2(new_n209_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n676_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n687_), .A2(new_n653_), .A3(new_n688_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n207_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n655_), .A2(KEYINPUT104), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n655_), .A2(KEYINPUT104), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n675_), .A2(new_n207_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n692_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(KEYINPUT46), .C1(new_n207_), .C2(new_n693_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1329gat));
  XNOR2_X1  g503(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n383_), .A2(new_n205_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n687_), .A2(new_n688_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n687_), .A2(KEYINPUT105), .A3(new_n688_), .A4(new_n706_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n383_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G43gat), .B1(new_n675_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AND4_X1   g512(.A1(new_n705_), .A2(new_n709_), .A3(new_n710_), .A4(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n705_), .B1(new_n715_), .B2(new_n710_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n687_), .A2(new_n472_), .A3(new_n688_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n556_), .A2(G50gat), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n718_), .A2(G50gat), .B1(new_n675_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT107), .ZN(G1331gat));
  NAND2_X1  g520(.A1(new_n623_), .A2(new_n624_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n614_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n628_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n634_), .A2(new_n637_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n583_), .A2(new_n608_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n331_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT108), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n331_), .A2(new_n730_), .A3(new_n727_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n642_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n727_), .A2(new_n648_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n641_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n738_), .A3(new_n697_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n697_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G64gat), .B1(new_n735_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1333gat));
  NOR2_X1   g542(.A1(new_n383_), .A2(G71gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n731_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G71gat), .B1(new_n735_), .B2(new_n383_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n732_), .A2(new_n752_), .A3(new_n472_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G78gat), .B1(new_n735_), .B2(new_n556_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1335gat));
  NAND2_X1  g555(.A1(new_n727_), .A2(new_n674_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT111), .ZN(new_n758_));
  INV_X1    g557(.A(G85gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n642_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n609_), .A2(new_n638_), .A3(new_n329_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n681_), .A2(new_n678_), .A3(new_n298_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n583_), .B2(new_n683_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n641_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n760_), .A2(new_n766_), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n758_), .A2(new_n499_), .A3(new_n653_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G92gat), .B1(new_n765_), .B2(new_n740_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1337gat));
  AND2_X1   g569(.A1(new_n711_), .A2(new_n230_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n764_), .A2(new_n711_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n758_), .A2(new_n771_), .B1(G99gat), .B2(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g573(.A1(new_n758_), .A2(new_n231_), .A3(new_n472_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n764_), .A2(new_n472_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n775_), .B(new_n781_), .C1(new_n779_), .C2(new_n778_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n589_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n586_), .A2(new_n587_), .A3(KEYINPUT55), .A4(new_n588_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n586_), .A2(new_n587_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT115), .B1(new_n789_), .B2(new_n590_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n791_), .B(new_n588_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n787_), .B(new_n788_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n599_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n796_), .A3(new_n599_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n620_), .A2(new_n618_), .A3(new_n629_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n615_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n723_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n725_), .A2(new_n601_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n795_), .A2(KEYINPUT58), .A3(new_n797_), .A4(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n789_), .A2(new_n590_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n791_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n789_), .A2(KEYINPUT115), .A3(new_n590_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n787_), .A2(new_n788_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n598_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n802_), .B1(new_n811_), .B2(new_n796_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n797_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n805_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n801_), .B1(new_n794_), .B2(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT58), .A4(new_n797_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n804_), .A2(new_n298_), .A3(new_n814_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n796_), .B1(new_n811_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n794_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n821_));
  INV_X1    g620(.A(new_n601_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n638_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n726_), .A2(new_n824_), .A3(new_n601_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n820_), .A2(new_n821_), .A3(new_n823_), .A4(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n602_), .A2(new_n725_), .A3(new_n800_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n647_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n818_), .B1(KEYINPUT57), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n819_), .B1(new_n793_), .B2(new_n599_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n823_), .B(new_n825_), .C1(new_n830_), .C2(KEYINPUT56), .ZN(new_n831_));
  INV_X1    g630(.A(new_n821_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n827_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n646_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n329_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT113), .B1(new_n329_), .B2(new_n726_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n638_), .A2(new_n840_), .A3(new_n328_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n608_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n683_), .B2(new_n842_), .ZN(new_n843_));
  AND4_X1   g642(.A1(new_n838_), .A2(new_n842_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n837_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n383_), .A2(new_n472_), .A3(new_n641_), .A4(new_n653_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n834_), .A2(new_n835_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n818_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n845_), .B1(new_n853_), .B2(new_n329_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT59), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n850_), .A2(new_n856_), .A3(new_n726_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G113gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n847_), .A2(new_n849_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n638_), .A2(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1340gat));
  NAND3_X1  g660(.A1(new_n850_), .A2(new_n856_), .A3(new_n609_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G120gat), .ZN(new_n863_));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(KEYINPUT60), .B2(new_n864_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n863_), .B1(new_n859_), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g666(.A(G127gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n328_), .B2(KEYINPUT118), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(KEYINPUT118), .B2(new_n868_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n850_), .A2(new_n856_), .A3(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n847_), .A2(new_n328_), .A3(new_n849_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(KEYINPUT119), .A3(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1342gat));
  AND2_X1   g677(.A1(new_n850_), .A2(new_n856_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT120), .B(G134gat), .Z(new_n880_));
  NOR2_X1   g679(.A1(new_n683_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n847_), .A2(new_n647_), .A3(new_n849_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n879_), .A2(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n711_), .A2(new_n556_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n854_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n697_), .A2(new_n641_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n726_), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n609_), .A3(new_n888_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g691(.A1(new_n887_), .A2(new_n328_), .A3(new_n888_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  NOR2_X1   g694(.A1(new_n646_), .A2(G162gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n887_), .A2(new_n888_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n888_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n854_), .A2(new_n683_), .A3(new_n886_), .A4(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(G162gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n897_), .B(KEYINPUT121), .C1(new_n900_), .C2(new_n899_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1347gat));
  NOR2_X1   g704(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n352_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n740_), .A2(new_n642_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n383_), .A2(new_n472_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n854_), .A2(new_n638_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n907_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n910_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n847_), .A2(new_n726_), .A3(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n906_), .B1(new_n913_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n912_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n906_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .A4(new_n907_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n911_), .A2(new_n344_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n854_), .A2(new_n910_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n609_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n328_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n355_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n336_), .B2(new_n927_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n847_), .A2(new_n914_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G190gat), .B1(new_n930_), .B2(new_n683_), .ZN(new_n931_));
  OR3_X1    g730(.A1(new_n646_), .A2(new_n515_), .A3(new_n514_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1351gat));
  NAND3_X1  g732(.A1(new_n887_), .A2(new_n726_), .A3(new_n908_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT124), .B1(new_n934_), .B2(new_n384_), .ZN(new_n935_));
  NOR4_X1   g734(.A1(new_n854_), .A2(new_n642_), .A3(new_n740_), .A4(new_n886_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n936_), .A2(new_n937_), .A3(G197gat), .A4(new_n726_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n934_), .A2(new_n384_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n935_), .A2(new_n938_), .A3(new_n939_), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n936_), .A2(new_n609_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n386_), .A2(KEYINPUT125), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT126), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n941_), .B(new_n943_), .ZN(G1353gat));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n328_), .B1(new_n945_), .B2(new_n302_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT127), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n936_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n945_), .A2(new_n302_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1354gat));
  NAND2_X1  g749(.A1(new_n887_), .A2(new_n908_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G218gat), .B1(new_n951_), .B2(new_n683_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n936_), .A2(new_n278_), .A3(new_n647_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1355gat));
endmodule


