//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT87), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(new_n203_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(KEYINPUT87), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n213_), .B(new_n214_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n215_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n208_), .B(new_n209_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n209_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n211_), .A2(new_n212_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n207_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n204_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n207_), .A2(KEYINPUT4), .A3(new_n226_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT99), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n228_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n233_), .A2(new_n234_), .B1(new_n236_), .B2(new_n230_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G85gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G57gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  NAND4_X1  g040(.A1(new_n229_), .A2(KEYINPUT99), .A3(new_n231_), .A4(new_n232_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT102), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n237_), .A2(KEYINPUT102), .A3(new_n241_), .A4(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n237_), .A2(new_n242_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G197gat), .A2(G204gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT91), .B(G197gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(G204gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(G211gat), .B(G218gat), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT21), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n256_), .A2(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(G197gat), .B2(G204gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n258_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(KEYINPUT21), .B2(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT79), .B(G183gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(G190gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT23), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n274_), .A2(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n270_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT85), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(KEYINPUT85), .ZN(new_n282_));
  AND2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n273_), .A2(KEYINPUT23), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n271_), .A2(KEYINPUT23), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI22_X1  g092(.A1(new_n288_), .A2(new_n291_), .B1(KEYINPUT24), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n283_), .A2(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n295_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n269_), .A2(KEYINPUT25), .ZN(new_n302_));
  OR2_X1    g101(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n269_), .A2(KEYINPUT80), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .A4(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n268_), .B1(new_n287_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n274_), .A2(new_n275_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n277_), .A2(new_n276_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n279_), .A3(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT96), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n300_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n297_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n293_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  OAI22_X1  g120(.A1(new_n288_), .A2(new_n291_), .B1(G183gat), .B2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n286_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n267_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n254_), .B1(new_n309_), .B2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n287_), .A2(new_n308_), .A3(new_n268_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n324_), .B2(new_n267_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n253_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT98), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n335_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT98), .ZN(new_n338_));
  INV_X1    g137(.A(new_n335_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n326_), .A2(new_n338_), .A3(new_n339_), .A4(new_n330_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n335_), .B(KEYINPUT103), .Z(new_n344_));
  NAND3_X1  g143(.A1(new_n327_), .A2(new_n254_), .A3(new_n329_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n267_), .B1(KEYINPUT100), .B2(new_n324_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT100), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n321_), .A2(new_n347_), .A3(new_n323_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n328_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n282_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n286_), .B1(new_n280_), .B2(KEYINPUT85), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n308_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n267_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n254_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT101), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n345_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI211_X1 g155(.A(KEYINPUT101), .B(new_n254_), .C1(new_n349_), .C2(new_n353_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n344_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT104), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n342_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n251_), .B(new_n343_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT30), .B1(new_n287_), .B2(new_n308_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n308_), .B(KEYINPUT30), .C1(new_n350_), .C2(new_n351_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT86), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G43gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G15gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n369_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n352_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT86), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n365_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n367_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT86), .B(new_n373_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT88), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n207_), .B(KEYINPUT31), .Z(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n226_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G22gat), .B(G50gat), .Z(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT93), .B1(G228gat), .B2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G78gat), .B(G106gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT94), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT93), .A2(G228gat), .A3(G233gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n267_), .B(new_n401_), .C1(new_n390_), .C2(new_n226_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT95), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n400_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n389_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n363_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n331_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n250_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n356_), .A2(new_n357_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n409_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n243_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n229_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n248_), .C1(new_n235_), .C2(new_n230_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n243_), .A2(new_n414_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n411_), .A2(new_n413_), .B1(new_n419_), .B2(new_n341_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n420_), .A2(new_n389_), .A3(new_n404_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n408_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G190gat), .B(G218gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G134gat), .B(G162gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT36), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G232gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(KEYINPUT35), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT10), .B(G99gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT64), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT65), .B(G85gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G92gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n436_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT6), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT7), .ZN(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n434_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n443_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT8), .ZN(new_n453_));
  XOR2_X1   g252(.A(G85gat), .B(G92gat), .Z(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT66), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n459_), .A3(new_n442_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n442_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n450_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n454_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT67), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n448_), .B(new_n449_), .C1(new_n466_), .C2(new_n442_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n465_), .B(new_n454_), .C1(new_n467_), .C2(new_n460_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(KEYINPUT8), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n455_), .B1(new_n469_), .B2(KEYINPUT68), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n464_), .A2(new_n471_), .A3(KEYINPUT8), .A4(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n445_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G29gat), .B(G36gat), .Z(new_n474_));
  XOR2_X1   g273(.A(G43gat), .B(G50gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n431_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n430_), .A2(KEYINPUT35), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n461_), .A2(new_n450_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n460_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n463_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT8), .B1(new_n481_), .B2(new_n465_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n468_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT68), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n455_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n472_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n444_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n476_), .B(KEYINPUT15), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n478_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n478_), .B1(new_n477_), .B2(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n426_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(KEYINPUT74), .B(new_n426_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n477_), .A2(new_n489_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n429_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n425_), .A2(KEYINPUT36), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n490_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n495_), .A2(new_n496_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n422_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n509_));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n510_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT69), .Z(new_n515_));
  AND3_X1   g314(.A1(new_n486_), .A2(new_n444_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n486_), .B2(new_n444_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n507_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT70), .B(new_n507_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n473_), .B2(new_n515_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n514_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n487_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n486_), .A2(new_n444_), .A3(new_n515_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n523_), .A2(new_n527_), .A3(new_n506_), .A4(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(new_n521_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n520_), .A2(new_n521_), .A3(new_n529_), .A4(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n535_), .B(new_n537_), .C1(KEYINPUT72), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT76), .B(G8gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT75), .B(G1gat), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G15gat), .B(G22gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n476_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(G229gat), .A3(G233gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n488_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n476_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G113gat), .B(G141gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n556_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT78), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT78), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n556_), .A2(new_n560_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n544_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n515_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n554_), .B(new_n580_), .Z(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT77), .Z(new_n584_));
  AND2_X1   g383(.A1(new_n581_), .A2(new_n514_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n581_), .A2(new_n514_), .ZN(new_n586_));
  NOR4_X1   g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n577_), .A4(new_n576_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n572_), .A2(KEYINPUT105), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n572_), .A2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT105), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n505_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n251_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n493_), .A2(KEYINPUT37), .A3(new_n502_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n503_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n588_), .ZN(new_n600_));
  NOR4_X1   g399(.A1(new_n422_), .A2(new_n571_), .A3(new_n544_), .A4(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n547_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n250_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  XNOR2_X1  g406(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n343_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n505_), .A2(new_n589_), .A3(new_n609_), .A4(new_n592_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G8gat), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n611_), .A2(KEYINPUT39), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(KEYINPUT39), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n546_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n608_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n616_), .B(new_n608_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1325gat));
  INV_X1    g419(.A(new_n389_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n371_), .B1(new_n593_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n601_), .A2(new_n371_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n601_), .A2(new_n626_), .A3(new_n405_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n593_), .A2(new_n405_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(G22gat), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT42), .B(new_n626_), .C1(new_n593_), .C2(new_n405_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  INV_X1    g433(.A(new_n599_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT108), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n599_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n636_), .B(new_n638_), .C1(new_n408_), .C2(new_n421_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n420_), .A2(new_n389_), .A3(new_n404_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n407_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n404_), .B1(new_n388_), .B2(new_n386_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n643_), .B2(new_n363_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n599_), .A2(KEYINPUT43), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n639_), .A2(KEYINPUT43), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n588_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n572_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n634_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n648_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n636_), .A2(new_n638_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n644_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n645_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n422_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n650_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n250_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n649_), .A2(KEYINPUT109), .A3(new_n250_), .A4(new_n656_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(G29gat), .A3(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n544_), .A2(new_n588_), .A3(new_n503_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n644_), .A2(new_n570_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G29gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n250_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n668_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n609_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n663_), .A2(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT45), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(KEYINPUT45), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n674_), .A2(new_n675_), .B1(KEYINPUT111), .B2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n649_), .A2(new_n609_), .A3(new_n656_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G36gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n676_), .A2(KEYINPUT111), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1329gat));
  NAND3_X1  g481(.A1(new_n649_), .A2(new_n621_), .A3(new_n656_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G43gat), .ZN(new_n684_));
  INV_X1    g483(.A(G43gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n663_), .A2(new_n685_), .A3(new_n621_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n663_), .B2(new_n405_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n649_), .A2(new_n656_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n405_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NAND3_X1  g491(.A1(new_n644_), .A2(new_n571_), .A3(new_n544_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n600_), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n250_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n543_), .A2(new_n647_), .A3(new_n570_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n505_), .A2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n250_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n695_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n698_), .B2(new_n609_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT48), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n701_), .A3(new_n609_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1333gat));
  NOR2_X1   g504(.A1(new_n389_), .A2(G71gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT112), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n694_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n698_), .A2(new_n621_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n698_), .B2(new_n405_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n694_), .A2(new_n716_), .A3(new_n405_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1335gat));
  NOR3_X1   g519(.A1(new_n693_), .A2(new_n588_), .A3(new_n503_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G85gat), .B1(new_n721_), .B2(new_n250_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n639_), .A2(KEYINPUT43), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n644_), .A2(new_n645_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n543_), .A2(new_n570_), .A3(new_n588_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n250_), .A2(new_n437_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n722_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  INV_X1    g528(.A(G92gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n721_), .A2(new_n730_), .A3(new_n609_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n727_), .A2(new_n609_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n730_), .ZN(G1337gat));
  AOI21_X1  g532(.A(new_n447_), .B1(new_n727_), .B2(new_n621_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n621_), .A2(new_n433_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n721_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n721_), .A2(new_n434_), .A3(new_n405_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n405_), .B(new_n726_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n434_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n725_), .A2(KEYINPUT114), .A3(new_n405_), .A4(new_n726_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT53), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n739_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n528_), .B1(new_n473_), .B2(new_n525_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n522_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n487_), .B2(new_n579_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n507_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT115), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n507_), .C1(new_n753_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n529_), .A2(KEYINPUT55), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n525_), .B1(new_n486_), .B2(new_n444_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n516_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n506_), .A4(new_n523_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n757_), .A2(new_n759_), .B1(new_n760_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n752_), .B1(new_n765_), .B2(new_n536_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n536_), .A2(new_n752_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT116), .B1(new_n765_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770_));
  INV_X1    g569(.A(new_n759_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n523_), .A2(new_n528_), .A3(new_n527_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n758_), .B1(new_n772_), .B2(new_n507_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n760_), .A2(new_n764_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n770_), .B(new_n767_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n766_), .A2(new_n769_), .A3(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n570_), .A2(new_n537_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n557_), .A2(new_n559_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n558_), .B1(new_n780_), .B2(KEYINPUT117), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(KEYINPUT117), .B2(new_n780_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n563_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n565_), .A2(new_n566_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n538_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n504_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n785_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n791_), .B2(new_n504_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n784_), .A2(new_n537_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n760_), .A2(new_n764_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n773_), .B2(new_n771_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n534_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n765_), .A2(new_n768_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n599_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI221_X1 g599(.A(new_n793_), .B1(KEYINPUT118), .B2(KEYINPUT58), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n789_), .A2(new_n792_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n647_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n543_), .A2(new_n599_), .A3(new_n571_), .A4(new_n588_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n609_), .A2(new_n251_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n641_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n570_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n807_), .B1(new_n803_), .B2(new_n647_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT59), .B1(new_n817_), .B2(new_n811_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n820_));
  AOI22_X1  g619(.A1(new_n786_), .A2(new_n788_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n588_), .B1(new_n821_), .B2(new_n792_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n812_), .B(new_n820_), .C1(new_n822_), .C2(new_n807_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n818_), .A2(new_n819_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n571_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n816_), .B1(new_n826_), .B2(new_n815_), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n823_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G120gat), .B1(new_n828_), .B2(new_n543_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G120gat), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n543_), .A2(KEYINPUT60), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n813_), .B2(new_n833_), .ZN(G1341gat));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n814_), .A2(new_n835_), .A3(new_n588_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n824_), .A2(new_n825_), .A3(new_n647_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(G1342gat));
  NAND2_X1  g637(.A1(new_n635_), .A2(G134gat), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n824_), .A2(new_n825_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT121), .B(new_n841_), .C1(new_n813_), .C2(new_n503_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n817_), .A2(new_n503_), .A3(new_n811_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G134gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT122), .B1(new_n840_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n818_), .A2(new_n819_), .A3(new_n823_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(G134gat), .A4(new_n635_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n842_), .A2(new_n845_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n847_), .A2(new_n853_), .ZN(G1343gat));
  NAND3_X1  g653(.A1(new_n809_), .A2(new_n642_), .A3(new_n810_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT123), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n817_), .A2(new_n406_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n810_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n571_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n211_), .ZN(G1344gat));
  AOI21_X1  g660(.A(new_n543_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n212_), .ZN(G1345gat));
  AOI21_X1  g662(.A(new_n647_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  NAND2_X1  g665(.A1(new_n856_), .A2(new_n859_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n867_), .A2(G162gat), .A3(new_n652_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n504_), .ZN(new_n869_));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(KEYINPUT124), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n503_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G162gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n868_), .B1(new_n871_), .B2(new_n874_), .ZN(G1347gat));
  NAND2_X1  g674(.A1(new_n609_), .A2(new_n251_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n817_), .A2(new_n407_), .A3(new_n876_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT125), .Z(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n284_), .A3(new_n570_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n570_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G169gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n285_), .A3(new_n544_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n877_), .A2(new_n544_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n285_), .B2(new_n886_), .ZN(G1349gat));
  AOI21_X1  g686(.A(new_n269_), .B1(new_n877_), .B2(new_n588_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n647_), .A2(new_n315_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n878_), .B2(new_n889_), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n878_), .A2(new_n300_), .A3(new_n504_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n877_), .B(KEYINPUT125), .ZN(new_n892_));
  OAI21_X1  g691(.A(G190gat), .B1(new_n892_), .B2(new_n599_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n817_), .A2(new_n406_), .A3(new_n876_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n570_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n544_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n588_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT63), .B(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n895_), .A2(new_n588_), .A3(new_n903_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n901_), .A2(new_n902_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n895_), .A2(new_n908_), .A3(new_n504_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n895_), .A2(new_n635_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1355gat));
endmodule


