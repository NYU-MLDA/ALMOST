//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n204_), .A2(new_n205_), .A3(G43gat), .ZN(new_n206_));
  INV_X1    g005(.A(G43gat), .ZN(new_n207_));
  INV_X1    g006(.A(G29gat), .ZN(new_n208_));
  INV_X1    g007(.A(G36gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n207_), .B1(new_n210_), .B2(new_n203_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n202_), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(G43gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n207_), .A3(new_n203_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(G50gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n212_), .A2(KEYINPUT15), .A3(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT15), .B1(new_n212_), .B2(new_n215_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219_));
  INV_X1    g018(.A(G1gat), .ZN(new_n220_));
  INV_X1    g019(.A(G8gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G1gat), .B(G8gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT76), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n212_), .A2(new_n215_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT75), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n225_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(G229gat), .A3(G233gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G169gat), .B(G197gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT77), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G113gat), .ZN(new_n238_));
  INV_X1    g037(.A(G141gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n232_), .A2(new_n234_), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT35), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n229_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  XOR2_X1   g051(.A(G85gat), .B(G92gat), .Z(new_n253_));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254_));
  AND3_X1   g053(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT65), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G99gat), .A2(G106gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n265_));
  NOR2_X1   g064(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI22_X1  g066(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n253_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT8), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT8), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n255_), .A2(new_n256_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n253_), .C1(new_n269_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT10), .B(G99gat), .Z(new_n277_));
  INV_X1    g076(.A(G106gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n253_), .A2(KEYINPUT9), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT9), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(G85gat), .A3(G92gat), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .A4(new_n273_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n252_), .B1(new_n276_), .B2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n257_), .A2(new_n262_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n272_), .B1(new_n285_), .B2(new_n253_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n253_), .A2(new_n272_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n267_), .A2(new_n268_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n273_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n252_), .B(new_n283_), .C1(new_n286_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n251_), .B1(new_n284_), .B2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT69), .B1(new_n247_), .B2(new_n248_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n283_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n295_), .B2(new_n218_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n250_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n283_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT66), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n229_), .B1(new_n300_), .B2(new_n290_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n301_), .A2(new_n249_), .A3(new_n296_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT70), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G190gat), .B(G218gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G134gat), .ZN(new_n305_));
  INV_X1    g104(.A(G162gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT36), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n292_), .A2(new_n250_), .A3(new_n297_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n249_), .B1(new_n301_), .B2(new_n296_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT37), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n307_), .A2(new_n308_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n317_), .A2(new_n318_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n309_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT37), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT13), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G57gat), .B(G64gat), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT11), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(KEYINPUT11), .ZN(new_n331_));
  XOR2_X1   g130(.A(G71gat), .B(G78gat), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n300_), .A2(new_n290_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n284_), .B2(new_n291_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G230gat), .A2(G233gat), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n295_), .A2(new_n338_), .A3(new_n335_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .A4(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n300_), .A2(new_n290_), .A3(new_n336_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n336_), .B1(new_n300_), .B2(new_n290_), .ZN(new_n346_));
  OAI211_X1 g145(.A(G230gat), .B(G233gat), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT67), .B(G204gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G120gat), .B(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT5), .B(G176gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(new_n347_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT68), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n344_), .A2(new_n347_), .A3(new_n355_), .A4(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n352_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n328_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  AOI211_X1 g159(.A(KEYINPUT13), .B(new_n358_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G231gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT72), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n225_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n225_), .A2(new_n364_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n335_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n336_), .A3(new_n366_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT16), .B(G183gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G211gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G155gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT17), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n368_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(KEYINPUT17), .A3(new_n376_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n327_), .A2(new_n362_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n244_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G127gat), .A2(G134gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G127gat), .A2(G134gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(G113gat), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G127gat), .ZN(new_n392_));
  INV_X1    g191(.A(G134gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G113gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n388_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n391_), .A2(new_n396_), .A3(G120gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(G120gat), .B1(new_n391_), .B2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n387_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n396_), .ZN(new_n400_));
  INV_X1    g199(.A(G120gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n396_), .A3(G120gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT83), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n399_), .A2(new_n404_), .A3(KEYINPUT31), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT31), .B1(new_n399_), .B2(new_n404_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT82), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT30), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT22), .B(G169gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n416_));
  INV_X1    g215(.A(G176gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n416_), .B2(KEYINPUT22), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G169gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT80), .ZN(new_n422_));
  OR2_X1    g221(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n423_));
  NAND2_X1  g222(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(G183gat), .B2(G190gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n418_), .A2(new_n436_), .A3(new_n420_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439_));
  NOR3_X1   g238(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n451_));
  AND2_X1   g250(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n423_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n427_), .A2(new_n429_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n446_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n438_), .A2(new_n439_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n439_), .B1(new_n438_), .B2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n414_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n458_), .A3(new_n413_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n411_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n464_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n471_), .A2(new_n409_), .A3(new_n410_), .A4(new_n466_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT1), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n479_), .B2(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(G148gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n239_), .A2(new_n482_), .A3(KEYINPUT84), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(G141gat), .B2(G148gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n480_), .A2(KEYINPUT85), .A3(new_n481_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G155gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n306_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n475_), .A3(new_n474_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n477_), .A2(KEYINPUT1), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n490_), .A3(new_n481_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(G141gat), .B2(G148gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n239_), .A3(new_n482_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT2), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n481_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n479_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n487_), .A2(new_n494_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT29), .ZN(new_n506_));
  INV_X1    g305(.A(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(G228gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(G228gat), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G211gat), .ZN(new_n514_));
  INV_X1    g313(.A(G218gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G211gat), .A2(G218gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT21), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G197gat), .B(G204gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT21), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(new_n522_), .A3(new_n517_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n518_), .A2(new_n520_), .A3(KEYINPUT21), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT89), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n525_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND4_X1   g329(.A1(new_n506_), .A2(new_n513_), .A3(new_n527_), .A4(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n513_), .B1(new_n506_), .B2(new_n528_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n531_), .A2(G78gat), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G78gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n506_), .A2(new_n528_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n512_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n506_), .A2(new_n513_), .A3(new_n527_), .A4(new_n530_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n278_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540_));
  OAI21_X1  g339(.A(G78gat), .B1(new_n531_), .B2(new_n532_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(G106gat), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n505_), .A2(KEYINPUT29), .ZN(new_n545_));
  XOR2_X1   g344(.A(G22gat), .B(G50gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT28), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n545_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .A4(new_n548_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n438_), .A2(new_n457_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n527_), .A2(new_n530_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT90), .B1(new_n452_), .B2(new_n451_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n558_));
  INV_X1    g357(.A(G190gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n561_));
  NAND2_X1  g360(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n449_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n430_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n445_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n415_), .A2(new_n417_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n442_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n433_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n528_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G226gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT19), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n554_), .A2(new_n555_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n574_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n566_), .A2(new_n570_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n553_), .B1(new_n579_), .B2(new_n526_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G8gat), .B(G36gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(G64gat), .B(G92gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n575_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n556_), .A2(new_n578_), .A3(new_n571_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n557_), .A2(new_n563_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n450_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n432_), .A3(new_n446_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n569_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n443_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n596_), .A3(KEYINPUT94), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n597_), .A3(new_n526_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT20), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n577_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n588_), .B1(new_n603_), .B2(new_n574_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT27), .B(new_n587_), .C1(new_n604_), .C2(new_n586_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT27), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n575_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n586_), .B1(new_n575_), .B2(new_n581_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n399_), .A2(new_n404_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n505_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n492_), .B(KEYINPUT85), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n397_), .A2(new_n398_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n504_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G225gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT92), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n613_), .A2(new_n504_), .B1(new_n404_), .B2(new_n399_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n614_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n505_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT4), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT4), .B1(new_n611_), .B2(new_n505_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n620_), .B1(new_n627_), .B2(new_n617_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT0), .B(G57gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G85gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(G1gat), .B(G29gat), .Z(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n612_), .A2(new_n615_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n625_), .B1(new_n635_), .B2(KEYINPUT4), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n619_), .B(new_n633_), .C1(new_n636_), .C2(new_n618_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n619_), .B1(new_n636_), .B2(new_n618_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n632_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n552_), .A2(new_n610_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n550_), .A2(new_n551_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n586_), .A2(KEYINPUT32), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n604_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n575_), .A2(new_n581_), .A3(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n645_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n576_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n578_), .B1(new_n649_), .B2(new_n602_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT96), .B(new_n648_), .C1(new_n650_), .C2(new_n588_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n641_), .A2(new_n646_), .A3(new_n647_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT93), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n637_), .B(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n607_), .A2(new_n608_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n627_), .A2(new_n618_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n632_), .C1(new_n618_), .C2(new_n635_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n643_), .B1(new_n652_), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n473_), .B1(new_n642_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n634_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n469_), .A2(new_n472_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n663_), .A2(new_n551_), .A3(new_n550_), .A4(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n665_), .B2(new_n610_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n610_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n473_), .A2(new_n641_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n552_), .A4(KEYINPUT98), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n661_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n386_), .B(new_n671_), .C1(new_n385_), .C2(new_n384_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT99), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(KEYINPUT99), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n675_), .A2(G1gat), .A3(new_n663_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT38), .Z(new_n677_));
  NOR2_X1   g476(.A1(new_n362_), .A2(new_n244_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n315_), .A2(new_n319_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT100), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT100), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n383_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n671_), .A2(new_n678_), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G1gat), .B1(new_n684_), .B2(new_n663_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n685_), .ZN(G1324gat));
  OAI21_X1  g485(.A(G8gat), .B1(new_n684_), .B2(new_n667_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT39), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n673_), .A2(new_n221_), .A3(new_n610_), .A4(new_n674_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT101), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT101), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  NOR3_X1   g493(.A1(new_n675_), .A2(G15gat), .A3(new_n473_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G15gat), .B1(new_n684_), .B2(new_n473_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT41), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT102), .Z(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n684_), .B2(new_n552_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n552_), .A2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n675_), .B2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n661_), .A2(KEYINPUT103), .A3(new_n670_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT103), .B1(new_n661_), .B2(new_n670_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n327_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n320_), .A2(new_n324_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT71), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(KEYINPUT43), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT104), .B1(new_n671_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n671_), .A2(KEYINPUT104), .A3(new_n713_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n678_), .B(new_n383_), .C1(new_n708_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n671_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n661_), .A2(new_n670_), .A3(KEYINPUT103), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n327_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT43), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n671_), .A2(KEYINPUT104), .A3(new_n713_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n714_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT44), .A3(new_n678_), .A4(new_n383_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n641_), .A3(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT105), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT105), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(G29gat), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n682_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n382_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n671_), .A3(new_n678_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n208_), .A3(new_n641_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n733_), .A2(new_n742_), .ZN(G1328gat));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT107), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n720_), .A2(new_n610_), .A3(new_n729_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G36gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(KEYINPUT107), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n738_), .A2(new_n209_), .A3(new_n610_), .A4(new_n739_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AND4_X1   g551(.A1(new_n745_), .A2(new_n747_), .A3(new_n748_), .A4(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n746_), .B2(G36gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n745_), .B1(new_n754_), .B2(new_n748_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1329gat));
  NAND4_X1  g555(.A1(new_n720_), .A2(G43gat), .A3(new_n664_), .A4(new_n729_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n207_), .B1(new_n740_), .B2(new_n473_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g559(.A1(new_n741_), .A2(new_n202_), .A3(new_n643_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n720_), .A2(new_n643_), .A3(new_n729_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n202_), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n241_), .A2(new_n243_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n661_), .B2(new_n670_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(new_n362_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n683_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n663_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n712_), .A2(new_n362_), .A3(new_n382_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT108), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n765_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(G57gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n772_), .B2(new_n663_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT109), .Z(G1332gat));
  OAI21_X1  g573(.A(G64gat), .B1(new_n767_), .B2(new_n667_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT48), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n667_), .A2(G64gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n771_), .B2(new_n777_), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n767_), .B2(new_n473_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT49), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n473_), .A2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n771_), .B2(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n767_), .B2(new_n552_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT110), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n643_), .A2(new_n534_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n786_), .B(new_n787_), .C1(new_n771_), .C2(new_n788_), .ZN(G1335gat));
  AND2_X1   g588(.A1(new_n766_), .A2(new_n735_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n641_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n362_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(new_n382_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n728_), .A2(new_n244_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n764_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n797_), .B2(new_n793_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n641_), .A2(G85gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n791_), .B1(new_n799_), .B2(new_n800_), .ZN(G1336gat));
  AOI21_X1  g600(.A(G92gat), .B1(new_n790_), .B2(new_n610_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n610_), .A2(G92gat), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT112), .Z(new_n804_));
  AOI21_X1  g603(.A(new_n802_), .B1(new_n799_), .B2(new_n804_), .ZN(G1337gat));
  NAND2_X1  g604(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G99gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n799_), .B2(new_n664_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n664_), .A2(new_n277_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n790_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n794_), .B(new_n795_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G99gat), .B1(new_n814_), .B2(new_n473_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n806_), .A3(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(G1338gat));
  OAI21_X1  g616(.A(G106gat), .B1(new_n794_), .B2(new_n552_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n790_), .A2(new_n278_), .A3(new_n643_), .ZN(new_n822_));
  OAI211_X1 g621(.A(G106gat), .B(new_n819_), .C1(new_n794_), .C2(new_n552_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n346_), .A2(new_n342_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n341_), .B1(new_n827_), .B2(new_n339_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n344_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n827_), .A2(KEYINPUT55), .A3(new_n341_), .A4(new_n339_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n352_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n357_), .B1(new_n833_), .B2(KEYINPUT56), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n244_), .B1(new_n833_), .B2(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n357_), .A2(new_n359_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n233_), .A2(new_n228_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n227_), .A2(new_n231_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n240_), .B(new_n838_), .C1(new_n839_), .C2(new_n228_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n243_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n835_), .A2(new_n836_), .B1(new_n837_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n826_), .B1(new_n843_), .B2(new_n682_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n842_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n836_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n834_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n734_), .A3(KEYINPUT57), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n832_), .B2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n357_), .C1(new_n849_), .C2(new_n832_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n852_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n327_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n844_), .A2(new_n848_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n383_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n764_), .A2(new_n383_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n327_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n327_), .C2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n244_), .A2(new_n382_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n837_), .A2(KEYINPUT13), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n357_), .A2(new_n328_), .A3(new_n359_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n712_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n868_), .A2(new_n712_), .A3(KEYINPUT115), .A4(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n864_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n864_), .B2(new_n874_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n857_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n610_), .A2(new_n663_), .A3(new_n473_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n552_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G113gat), .B1(new_n881_), .B2(new_n764_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(G113gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n864_), .A2(new_n874_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT117), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n864_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n643_), .B1(new_n889_), .B2(new_n857_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n885_), .B1(new_n890_), .B2(new_n879_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AND4_X1   g692(.A1(new_n552_), .A2(new_n878_), .A3(new_n879_), .A4(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n880_), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n890_), .A2(new_n879_), .A3(new_n893_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n884_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G113gat), .B1(new_n244_), .B2(new_n883_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n882_), .B1(new_n900_), .B2(new_n901_), .ZN(G1340gat));
  OAI21_X1  g701(.A(new_n401_), .B1(new_n792_), .B2(KEYINPUT60), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n881_), .B(new_n903_), .C1(KEYINPUT60), .C2(new_n401_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n891_), .A2(new_n894_), .A3(new_n792_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n401_), .ZN(G1341gat));
  NAND3_X1  g705(.A1(new_n881_), .A2(new_n392_), .A3(new_n382_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n383_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n392_), .ZN(G1342gat));
  NAND3_X1  g708(.A1(new_n881_), .A2(new_n393_), .A3(new_n682_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n712_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n393_), .ZN(G1343gat));
  AOI21_X1  g711(.A(new_n664_), .B1(new_n889_), .B2(new_n857_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n552_), .A2(new_n610_), .A3(new_n663_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n244_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT122), .B(G141gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1344gat));
  NOR2_X1   g717(.A1(new_n915_), .A2(new_n792_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n482_), .ZN(G1345gat));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n913_), .A2(new_n921_), .A3(new_n382_), .A4(new_n914_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n878_), .A2(new_n473_), .A3(new_n382_), .A4(new_n914_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT123), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n922_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n488_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n924_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT61), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n922_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(G155gat), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n932_), .ZN(G1346gat));
  NOR3_X1   g732(.A1(new_n915_), .A2(new_n306_), .A3(new_n712_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n913_), .A2(new_n682_), .A3(new_n914_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n306_), .B2(new_n935_), .ZN(G1347gat));
  NAND4_X1  g735(.A1(new_n878_), .A2(new_n552_), .A3(new_n610_), .A4(new_n668_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n764_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(G169gat), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n938_), .A2(new_n764_), .A3(new_n415_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n942_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n939_), .A2(G169gat), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n943_), .A2(new_n944_), .A3(new_n947_), .ZN(G1348gat));
  NOR2_X1   g747(.A1(new_n937_), .A2(new_n792_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(new_n417_), .ZN(G1349gat));
  NOR2_X1   g749(.A1(new_n937_), .A2(new_n383_), .ZN(new_n951_));
  MUX2_X1   g750(.A(G183gat), .B(new_n450_), .S(new_n951_), .Z(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n937_), .B2(new_n712_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n682_), .A2(new_n591_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n937_), .B2(new_n954_), .ZN(G1351gat));
  AND3_X1   g754(.A1(new_n878_), .A2(new_n610_), .A3(new_n473_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n552_), .A2(new_n641_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n764_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n956_), .A2(new_n957_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n792_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(G204gat), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n963_), .A2(G204gat), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n962_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n966_), .B1(new_n962_), .B2(new_n964_), .ZN(G1353gat));
  AOI21_X1  g766(.A(new_n383_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT126), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  OR2_X1    g771(.A1(new_n970_), .A2(new_n971_), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n958_), .A2(new_n968_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n956_), .A2(new_n957_), .A3(new_n968_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n972_), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n958_), .B2(new_n682_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n961_), .A2(new_n515_), .A3(new_n712_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1355gat));
endmodule


