//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G183gat), .B(G211gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT17), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(KEYINPUT17), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT14), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G1gat), .ZN(new_n213_));
  INV_X1    g012(.A(G8gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n210_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .A4(new_n215_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G64gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G57gat), .ZN(new_n223_));
  INV_X1    g022(.A(G57gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G64gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n227_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT11), .B1(new_n223_), .B2(new_n225_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G78gat), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n233_), .A2(KEYINPUT67), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n228_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n233_), .B2(new_n234_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n228_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n221_), .B(new_n241_), .ZN(new_n242_));
  MUX2_X1   g041(.A(new_n207_), .B(new_n208_), .S(new_n242_), .Z(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT79), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G43gat), .B(G50gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n247_), .B(new_n249_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260_));
  AND2_X1   g059(.A1(G85gat), .A2(G92gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G85gat), .A2(G92gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G85gat), .ZN(new_n264_));
  INV_X1    g063(.A(G92gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT66), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G99gat), .A2(G106gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT7), .ZN(new_n274_));
  INV_X1    g073(.A(G99gat), .ZN(new_n275_));
  INV_X1    g074(.A(G106gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n279_));
  AND4_X1   g078(.A1(new_n273_), .A2(new_n277_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT8), .B1(new_n270_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n266_), .A2(new_n267_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT65), .B1(new_n283_), .B2(new_n260_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT8), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n277_), .A2(new_n273_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .A4(new_n268_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n281_), .A2(new_n282_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT9), .B1(new_n261_), .B2(new_n262_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT9), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n267_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT10), .B(G99gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n273_), .B(new_n278_), .C1(new_n294_), .C2(G106gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n290_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n288_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n282_), .B1(new_n281_), .B2(new_n287_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n259_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT34), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT72), .Z(new_n305_));
  NOR2_X1   g104(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n281_), .A2(new_n287_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n256_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n301_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n301_), .B2(new_n308_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(KEYINPUT36), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n246_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n301_), .A2(new_n308_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n305_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n301_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n246_), .A3(new_n315_), .A4(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n314_), .B(KEYINPUT36), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n316_), .A2(new_n322_), .B1(new_n311_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n324_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n319_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT74), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n330_), .B2(new_n321_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT37), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT76), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT76), .B1(new_n309_), .B2(new_n310_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n323_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(new_n321_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n245_), .B1(new_n334_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n281_), .A2(new_n287_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n298_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n239_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT68), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n307_), .A2(new_n241_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n347_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G230gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n345_), .A2(new_n346_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n307_), .A2(new_n241_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n307_), .B2(new_n241_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(new_n353_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G120gat), .B(G148gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT5), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G176gat), .B(G204gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n355_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n361_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n349_), .B1(new_n307_), .B2(new_n241_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(new_n359_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n353_), .B1(new_n373_), .B2(new_n350_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n355_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT70), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT13), .B1(new_n370_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(KEYINPUT70), .A3(new_n376_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT13), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n378_), .A2(KEYINPUT71), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT71), .B1(new_n378_), .B2(new_n382_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OR3_X1    g184(.A1(new_n342_), .A2(new_n385_), .A3(KEYINPUT80), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT80), .B1(new_n342_), .B2(new_n385_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  INV_X1    g187(.A(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(G15gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n390_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT25), .B(G183gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G169gat), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT24), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n398_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT23), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(KEYINPUT24), .B2(new_n405_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n398_), .B(KEYINPUT84), .C1(new_n402_), .C2(new_n406_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT22), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(G169gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n404_), .B1(new_n420_), .B2(KEYINPUT85), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT22), .B(G169gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(KEYINPUT85), .B2(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n414_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n401_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(new_n399_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n418_), .A2(new_n431_), .A3(KEYINPUT30), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT30), .B1(new_n418_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n395_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n418_), .A2(new_n431_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n394_), .A3(new_n432_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G127gat), .B(G134gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G113gat), .B(G120gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT31), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT86), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n435_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G204gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G197gat), .ZN(new_n455_));
  INV_X1    g254(.A(G197gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G204gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT21), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n456_), .B2(G204gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT21), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n458_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n455_), .A2(new_n457_), .A3(KEYINPUT94), .A4(KEYINPUT21), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n453_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI211_X1 g266(.A(KEYINPUT95), .B(new_n453_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n459_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G155gat), .A2(G162gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT88), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(G141gat), .ZN(new_n478_));
  INV_X1    g277(.A(G148gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .A4(KEYINPUT87), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n481_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT3), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n474_), .B1(new_n476_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n473_), .B1(new_n471_), .B2(KEYINPUT1), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(KEYINPUT1), .B2(new_n473_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G141gat), .B(G148gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n470_), .B1(new_n491_), .B2(KEYINPUT29), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n451_), .B1(new_n469_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n469_), .A2(new_n492_), .A3(new_n451_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G78gat), .B(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n495_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n498_), .B1(new_n499_), .B2(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(KEYINPUT96), .ZN(new_n502_));
  XOR2_X1   g301(.A(G22gat), .B(G50gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n486_), .A2(new_n507_), .A3(new_n490_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT89), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n486_), .A2(new_n511_), .A3(new_n507_), .A4(new_n490_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT91), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n505_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n501_), .A2(new_n502_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n519_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n500_), .B(new_n497_), .C1(new_n522_), .C2(KEYINPUT96), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n442_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n486_), .A2(new_n490_), .A3(new_n442_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G225gat), .A2(G233gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT100), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n526_), .A2(KEYINPUT4), .A3(new_n527_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n526_), .B2(KEYINPUT4), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT0), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G57gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n535_), .A2(KEYINPUT0), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(KEYINPUT0), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n224_), .A3(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n537_), .A2(new_n540_), .A3(G85gat), .ZN(new_n541_));
  AOI21_X1  g340(.A(G85gat), .B1(new_n537_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n545_), .B(new_n531_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n524_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT20), .ZN(new_n549_));
  INV_X1    g348(.A(new_n406_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n550_), .A2(new_n428_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n415_), .B1(new_n551_), .B2(KEYINPUT84), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n430_), .B1(new_n552_), .B2(new_n409_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n469_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n459_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n465_), .A2(new_n466_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n464_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n461_), .A2(KEYINPUT21), .B1(new_n455_), .B2(new_n457_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n452_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT95), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n555_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n400_), .A2(KEYINPUT98), .A3(new_n401_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n427_), .B2(new_n399_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n562_), .A2(new_n564_), .B1(new_n404_), .B2(new_n422_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n414_), .B2(new_n425_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n414_), .A2(new_n566_), .A3(new_n425_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n550_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n416_), .A2(new_n398_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n561_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n549_), .B1(new_n554_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G226gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT19), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n576_), .B(KEYINPUT97), .Z(new_n579_));
  INV_X1    g378(.A(new_n572_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT20), .B1(new_n580_), .B2(new_n561_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n436_), .A2(new_n469_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G8gat), .B(G36gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT18), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G64gat), .B(G92gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(KEYINPUT27), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n549_), .B1(new_n469_), .B2(new_n572_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n561_), .A2(new_n553_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n579_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n587_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n549_), .B(new_n576_), .C1(new_n554_), .C2(new_n573_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n592_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n588_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT27), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n589_), .A2(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n548_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(KEYINPUT32), .A3(new_n587_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n587_), .A2(KEYINPUT32), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n578_), .A2(new_n583_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n547_), .A3(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n532_), .A2(new_n533_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(KEYINPUT33), .A3(new_n531_), .A4(new_n545_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n543_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n543_), .B2(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n530_), .B1(new_n526_), .B2(KEYINPUT4), .ZN(new_n614_));
  OAI22_X1  g413(.A1(new_n612_), .A2(new_n613_), .B1(new_n532_), .B2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n599_), .A2(new_n588_), .A3(new_n609_), .A4(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n546_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n546_), .B2(new_n618_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n607_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n524_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n448_), .B1(new_n603_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n600_), .A2(new_n601_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n447_), .A2(new_n547_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n596_), .A2(KEYINPUT27), .A3(new_n588_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n524_), .A2(new_n625_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n602_), .A2(KEYINPUT103), .A3(new_n524_), .A4(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n624_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT81), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n219_), .B2(new_n253_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n256_), .A2(KEYINPUT81), .A3(new_n217_), .A4(new_n218_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n255_), .A2(new_n258_), .A3(new_n219_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT82), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT82), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n637_), .A2(new_n642_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n219_), .A2(new_n253_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n637_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n638_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n641_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G113gat), .B(G141gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G169gat), .B(G197gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n648_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n633_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n386_), .A2(new_n387_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n213_), .A3(new_n547_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n378_), .A2(new_n382_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n653_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n633_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n337_), .A2(new_n338_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n245_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n547_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(new_n667_), .ZN(G1324gat));
  INV_X1    g467(.A(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n602_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n214_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n657_), .A2(new_n214_), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1325gat));
  AOI21_X1  g476(.A(new_n392_), .B1(new_n669_), .B2(new_n448_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n392_), .A3(new_n448_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT105), .ZN(G1326gat));
  AND2_X1   g481(.A1(new_n524_), .A2(KEYINPUT106), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n524_), .A2(KEYINPUT106), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n665_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT42), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n686_), .A2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n656_), .B2(new_n689_), .ZN(G1327gat));
  INV_X1    g489(.A(new_n663_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n244_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n662_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n547_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n326_), .A2(new_n333_), .B1(new_n663_), .B2(new_n339_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n624_), .B2(new_n632_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT43), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n696_), .C1(new_n624_), .C2(new_n632_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n244_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n661_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(KEYINPUT44), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n705_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n547_), .A2(G29gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n695_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n602_), .A2(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n694_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n693_), .A2(KEYINPUT45), .A3(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n713_), .A2(KEYINPUT108), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n670_), .A3(new_n707_), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(KEYINPUT108), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT46), .ZN(G1329gat));
  NOR2_X1   g520(.A1(new_n447_), .A2(new_n389_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n707_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n389_), .B1(new_n693_), .B2(new_n447_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT109), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n723_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n726_), .B(new_n731_), .C1(new_n728_), .C2(new_n723_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n694_), .B2(new_n685_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n524_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n708_), .B2(new_n736_), .ZN(G1331gat));
  AOI22_X1  g536(.A1(new_n602_), .A2(new_n548_), .B1(new_n622_), .B2(new_n524_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n630_), .B(new_n631_), .C1(new_n738_), .C2(new_n448_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n660_), .A2(new_n653_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n341_), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n224_), .A3(new_n547_), .ZN(new_n742_));
  AND4_X1   g541(.A1(new_n664_), .A2(new_n385_), .A3(new_n739_), .A4(new_n654_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n547_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(new_n224_), .ZN(G1332gat));
  AOI21_X1  g544(.A(new_n222_), .B1(new_n743_), .B2(new_n670_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT48), .Z(new_n747_));
  NOR2_X1   g546(.A1(new_n602_), .A2(G64gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT110), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n741_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n743_), .B2(new_n448_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT49), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n741_), .A2(new_n752_), .A3(new_n448_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n743_), .B2(new_n685_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT50), .Z(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(new_n757_), .A3(new_n685_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1335gat));
  NAND4_X1  g560(.A1(new_n385_), .A2(new_n739_), .A3(new_n654_), .A4(new_n692_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n264_), .A3(new_n547_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n700_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n699_), .B1(new_n739_), .B2(new_n696_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n245_), .B(new_n740_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT112), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n701_), .A2(new_n770_), .A3(new_n740_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n666_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n765_), .B1(new_n772_), .B2(new_n264_), .ZN(G1336gat));
  NAND3_X1  g572(.A1(new_n764_), .A2(new_n265_), .A3(new_n670_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n602_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n265_), .ZN(G1337gat));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n768_), .A2(KEYINPUT112), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n701_), .B2(new_n740_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n448_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G99gat), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n447_), .A2(new_n294_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n764_), .A2(new_n785_), .B1(new_n777_), .B2(KEYINPUT51), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n780_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n447_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n780_), .B(new_n786_), .C1(new_n788_), .C2(new_n275_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n779_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n275_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n778_), .A3(new_n789_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n764_), .A2(new_n276_), .A3(new_n735_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n701_), .A2(new_n735_), .A3(new_n740_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G106gat), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n798_), .A3(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n797_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n797_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  NOR2_X1   g608(.A1(new_n670_), .A2(new_n735_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n547_), .A3(new_n448_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT75), .B1(new_n325_), .B2(KEYINPUT37), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n331_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n340_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n653_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n244_), .A4(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n341_), .A2(new_n819_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n244_), .A3(new_n816_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT54), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n653_), .A2(new_n376_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n361_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT12), .B1(new_n344_), .B2(new_n347_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n351_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT55), .A3(new_n353_), .A4(new_n358_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n828_), .A2(new_n358_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n826_), .B(new_n829_), .C1(new_n830_), .C2(new_n353_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n365_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n365_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n824_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n641_), .A2(new_n647_), .A3(new_n643_), .A4(new_n652_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n637_), .A2(new_n639_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT118), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n637_), .A2(new_n840_), .A3(new_n639_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n638_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n652_), .B1(new_n645_), .B2(new_n638_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n837_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n691_), .B1(new_n836_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n365_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n365_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n845_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT119), .A3(new_n376_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n367_), .B2(new_n845_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n850_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n834_), .A2(new_n835_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT58), .A3(new_n857_), .A4(new_n855_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n696_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n691_), .C1(new_n836_), .C2(new_n846_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n245_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n811_), .B1(new_n823_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n653_), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n811_), .C1(new_n823_), .C2(new_n865_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n823_), .A2(new_n865_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n811_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n866_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n868_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n653_), .A2(G113gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT121), .Z(new_n878_));
  AOI21_X1  g677(.A(new_n867_), .B1(new_n876_), .B2(new_n878_), .ZN(G1340gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n876_), .B2(new_n385_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(KEYINPUT60), .B2(new_n881_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n871_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n880_), .B1(new_n882_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n887_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n385_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n890_), .B(new_n868_), .C1(new_n873_), .C2(new_n875_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT123), .B(new_n889_), .C1(new_n891_), .C2(new_n881_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1341gat));
  AOI21_X1  g692(.A(G127gat), .B1(new_n866_), .B2(new_n244_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n244_), .A2(KEYINPUT124), .A3(G127gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(KEYINPUT124), .B2(G127gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n876_), .B2(new_n896_), .ZN(G1342gat));
  INV_X1    g696(.A(G134gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n866_), .A2(new_n898_), .A3(new_n663_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n876_), .A2(new_n696_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1343gat));
  NAND2_X1  g700(.A1(new_n735_), .A2(new_n447_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(new_n670_), .A3(new_n666_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n869_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n654_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n478_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n890_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n479_), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n245_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n904_), .B2(new_n814_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n691_), .A2(G162gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n904_), .B2(new_n913_), .ZN(G1347gat));
  NOR3_X1   g713(.A1(new_n602_), .A2(new_n547_), .A3(new_n447_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n686_), .A2(new_n653_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n403_), .B1(new_n869_), .B2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT62), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n602_), .B1(new_n823_), .B2(new_n865_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n920_), .A2(new_n626_), .A3(new_n686_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n422_), .A3(new_n653_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1348gat));
  INV_X1    g722(.A(new_n660_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G176gat), .B1(new_n921_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n869_), .A2(new_n524_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n385_), .A2(G176gat), .A3(new_n915_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n927_), .A2(new_n244_), .A3(new_n915_), .ZN(new_n930_));
  INV_X1    g729(.A(G183gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n245_), .A2(new_n396_), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n930_), .A2(new_n931_), .B1(new_n921_), .B2(new_n932_), .ZN(G1350gat));
  NAND2_X1  g732(.A1(new_n921_), .A2(new_n696_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G190gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n921_), .A2(new_n663_), .A3(new_n397_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n902_), .A2(new_n547_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n920_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n654_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n456_), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n890_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n454_), .ZN(G1353gat));
  INV_X1    g742(.A(new_n939_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n245_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(KEYINPUT125), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n946_), .A2(new_n947_), .A3(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(new_n949_), .B2(new_n946_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n947_), .B1(new_n946_), .B2(new_n949_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1354gat));
  XOR2_X1   g752(.A(KEYINPUT127), .B(G218gat), .Z(new_n954_));
  NOR3_X1   g753(.A1(new_n939_), .A2(new_n814_), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n944_), .A2(new_n663_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n954_), .ZN(G1355gat));
endmodule


