//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT72), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n212_));
  INV_X1    g011(.A(G57gat), .ZN(new_n213_));
  INV_X1    g012(.A(G64gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G57gat), .A2(G64gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(G78gat), .ZN(new_n221_));
  INV_X1    g020(.A(G78gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(new_n218_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n217_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n216_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G57gat), .A2(G64gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT11), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(G78gat), .B1(new_n219_), .B2(new_n220_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n212_), .A3(new_n216_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n211_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT16), .B(G183gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G211gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G155gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n241_), .B1(KEYINPUT17), .B2(new_n240_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G15gat), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT82), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT83), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT80), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261_));
  AOI21_X1  g060(.A(G176gat), .B1(new_n254_), .B2(new_n255_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n259_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  INV_X1    g064(.A(G190gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT23), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n264_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT25), .B(G183gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n266_), .B2(KEYINPUT26), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G190gat), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n274_), .B(new_n276_), .C1(new_n277_), .C2(new_n275_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n269_), .A2(KEYINPUT79), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT79), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(new_n268_), .A3(G183gat), .A4(G190gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n267_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n257_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n285_), .A2(KEYINPUT24), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n285_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n259_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n283_), .A2(new_n288_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n273_), .B1(new_n279_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n273_), .B(KEYINPUT81), .C1(new_n279_), .C2(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT30), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(KEYINPUT84), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(KEYINPUT84), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n253_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n298_), .B2(new_n253_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302_));
  INV_X1    g101(.A(G113gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G120gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT85), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n304_), .B(G120gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT31), .Z(new_n312_));
  AND2_X1   g111(.A1(new_n301_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n301_), .A2(new_n312_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(KEYINPUT2), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  OR3_X1    g118(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(KEYINPUT2), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G155gat), .ZN(new_n323_));
  INV_X1    g122(.A(G162gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT86), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(G155gat), .B2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT87), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G155gat), .A3(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  INV_X1    g135(.A(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n329_), .B(new_n336_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT88), .B1(new_n340_), .B2(new_n328_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n338_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n344_));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345_));
  AND3_X1   g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n335_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n348_), .A2(KEYINPUT29), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n348_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G197gat), .B(G204gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n353_), .A2(KEYINPUT21), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G197gat), .B(G204gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n354_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n357_), .A2(new_n358_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n354_), .B(new_n359_), .C1(new_n362_), .C2(new_n355_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n348_), .B2(KEYINPUT29), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  AOI211_X1 g167(.A(new_n368_), .B(new_n364_), .C1(new_n348_), .C2(KEYINPUT29), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G22gat), .B(G50gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT28), .Z(new_n371_));
  NOR3_X1   g170(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n364_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n335_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n343_), .A2(new_n345_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT89), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n368_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n365_), .A2(new_n366_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n373_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n352_), .B1(new_n372_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n371_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n383_), .A3(new_n373_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n351_), .A4(new_n350_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT18), .B(G64gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G92gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT98), .Z(new_n394_));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT19), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n283_), .A2(new_n271_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n259_), .A3(new_n258_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n277_), .A2(new_n274_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n289_), .A3(new_n286_), .A4(new_n270_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n364_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT97), .B1(new_n402_), .B2(KEYINPUT20), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n296_), .B2(new_n374_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n397_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n294_), .A2(new_n295_), .A3(new_n364_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n374_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(KEYINPUT20), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(new_n396_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n394_), .B1(new_n406_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n296_), .A2(new_n374_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n402_), .A2(KEYINPUT91), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n402_), .A2(KEYINPUT91), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n413_), .A2(new_n416_), .A3(new_n397_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n396_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n393_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n412_), .A2(KEYINPUT27), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n419_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n393_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n420_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT99), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n418_), .A2(new_n419_), .A3(new_n393_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n393_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT99), .B(new_n426_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n389_), .B(new_n421_), .C1(new_n427_), .C2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT93), .B1(new_n379_), .B2(new_n311_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n348_), .A2(new_n434_), .A3(new_n307_), .A4(new_n310_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n379_), .A2(new_n306_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n379_), .A2(new_n311_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT4), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n437_), .B2(KEYINPUT4), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT0), .B(G57gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G85gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(G1gat), .B(G29gat), .Z(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n438_), .B(new_n442_), .C1(KEYINPUT4), .C2(new_n437_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n439_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT100), .B1(new_n432_), .B2(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n451_), .A2(new_n450_), .A3(new_n439_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n443_), .A2(new_n440_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n439_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT100), .ZN(new_n460_));
  INV_X1    g259(.A(new_n421_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT99), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n464_), .B2(new_n430_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n459_), .A2(new_n460_), .A3(new_n389_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n454_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n437_), .A2(KEYINPUT4), .ZN(new_n469_));
  INV_X1    g268(.A(new_n442_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n440_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n433_), .A2(new_n435_), .A3(new_n440_), .A4(new_n436_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n448_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n468_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n475_), .B(KEYINPUT96), .C1(new_n443_), .C2(new_n440_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(KEYINPUT33), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n425_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT92), .B1(new_n424_), .B2(new_n420_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n480_), .B1(new_n478_), .B2(KEYINPUT33), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n450_), .B(new_n486_), .C1(new_n451_), .C2(new_n439_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n477_), .A2(new_n481_), .A3(new_n485_), .A4(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n422_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n406_), .B2(new_n411_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n490_), .B(new_n491_), .C1(new_n455_), .C2(new_n458_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n389_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n316_), .B1(new_n467_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n389_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n315_), .A2(new_n459_), .A3(new_n495_), .A4(new_n465_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n246_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(KEYINPUT10), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(KEYINPUT10), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT9), .ZN(new_n510_));
  INV_X1    g309(.A(G85gat), .ZN(new_n511_));
  INV_X1    g310(.A(G92gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(KEYINPUT9), .A3(new_n509_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n503_), .A2(new_n508_), .A3(new_n510_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n500_), .A3(new_n499_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n506_), .A3(new_n507_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n513_), .A2(new_n509_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n515_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n234_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n233_), .B(new_n515_), .C1(new_n523_), .C2(new_n522_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n498_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(KEYINPUT12), .A3(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n234_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT65), .B1(new_n532_), .B2(new_n498_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  INV_X1    g333(.A(new_n498_), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n534_), .B(new_n535_), .C1(new_n529_), .C2(new_n531_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n528_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G120gat), .B(G148gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n257_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n537_), .A2(KEYINPUT66), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT66), .B1(new_n537_), .B2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n528_), .B(new_n541_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT67), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT13), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT66), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n532_), .A2(new_n498_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n534_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n535_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT65), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n527_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n554_), .B2(new_n541_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n537_), .A2(KEYINPUT66), .A3(new_n542_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(KEYINPUT67), .A3(new_n541_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n546_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n548_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G29gat), .B(G36gat), .ZN(new_n566_));
  INV_X1    g365(.A(G43gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G50gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n566_), .B(G43gat), .ZN(new_n570_));
  INV_X1    g369(.A(G50gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT74), .ZN(new_n574_));
  INV_X1    g373(.A(new_n208_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT15), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n208_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT76), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n573_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n208_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n576_), .A3(KEYINPUT75), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n574_), .A2(KEYINPUT75), .A3(new_n575_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n583_), .B1(new_n589_), .B2(new_n581_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G169gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G197gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n590_), .B(new_n593_), .Z(new_n594_));
  NOR2_X1   g393(.A1(new_n565_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n497_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G134gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n324_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT36), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n573_), .A2(new_n524_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT70), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n578_), .A2(new_n524_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT68), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT34), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT71), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n603_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n606_), .A2(new_n608_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n600_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n599_), .A2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n613_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n596_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n203_), .A3(new_n453_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT38), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n616_), .A2(new_n620_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n596_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n459_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n465_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n204_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G8gat), .B1(new_n631_), .B2(new_n465_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(KEYINPUT39), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(KEYINPUT39), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g439(.A1(new_n625_), .A2(G15gat), .A3(new_n316_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n596_), .A2(new_n315_), .A3(new_n630_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(G15gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n642_), .A3(G15gat), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(KEYINPUT41), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT41), .B1(new_n645_), .B2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n641_), .B1(new_n647_), .B2(new_n648_), .ZN(G1326gat));
  NAND3_X1  g448(.A1(new_n596_), .A2(new_n389_), .A3(new_n630_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G22gat), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n625_), .A2(G22gat), .A3(new_n495_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT103), .ZN(G1327gat));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n623_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n494_), .A2(new_n496_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n623_), .B(KEYINPUT104), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n663_), .B1(new_n666_), .B2(KEYINPUT43), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n595_), .A2(new_n246_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT44), .B(new_n670_), .C1(new_n671_), .C2(new_n663_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n453_), .A3(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(KEYINPUT105), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(G29gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n630_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n668_), .ZN(new_n679_));
  INV_X1    g478(.A(G29gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n453_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n669_), .A2(new_n634_), .A3(new_n672_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n677_), .A2(new_n686_), .A3(new_n634_), .A4(new_n670_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT45), .Z(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(KEYINPUT106), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT46), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n688_), .B1(new_n684_), .B2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n691_), .B2(KEYINPUT46), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n683_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n693_), .A2(new_n695_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n693_), .B2(KEYINPUT106), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n698_), .B(KEYINPUT108), .C1(new_n699_), .C2(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n669_), .A2(new_n672_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G43gat), .B1(new_n702_), .B2(new_n316_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n679_), .A2(new_n567_), .A3(new_n315_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n702_), .B2(new_n495_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n679_), .A2(new_n571_), .A3(new_n389_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1331gat));
  XNOR2_X1  g508(.A(new_n590_), .B(new_n593_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n564_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n497_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n630_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n213_), .A3(new_n459_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n624_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n459_), .B1(new_n716_), .B2(KEYINPUT109), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(KEYINPUT109), .B2(new_n716_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n213_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n713_), .B2(new_n465_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n214_), .A3(new_n634_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n713_), .B2(new_n316_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n715_), .A2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n316_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n713_), .B2(new_n495_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n716_), .A2(new_n222_), .A3(new_n389_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  NAND2_X1  g530(.A1(new_n711_), .A2(new_n246_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n677_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n511_), .B1(new_n734_), .B2(new_n459_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT110), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n667_), .A2(new_n732_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n459_), .A2(new_n511_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(G1336gat));
  OAI21_X1  g538(.A(new_n512_), .B1(new_n734_), .B2(new_n465_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT111), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(G92gat), .A3(new_n634_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT112), .Z(G1337gat));
  NOR2_X1   g543(.A1(new_n501_), .A2(new_n502_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n734_), .A2(new_n745_), .A3(new_n316_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT113), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n500_), .B1(new_n737_), .B2(new_n315_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g549(.A(new_n499_), .B1(new_n737_), .B2(new_n389_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT52), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n734_), .A2(G106gat), .A3(new_n495_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT114), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n590_), .A2(new_n593_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n582_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n593_), .B1(new_n589_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT120), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n580_), .A2(new_n760_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n557_), .A2(new_n562_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT117), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n532_), .A2(new_n498_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n552_), .B2(KEYINPUT55), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n768_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n770_), .A2(KEYINPUT118), .A3(new_n772_), .A4(new_n774_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n542_), .A4(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n710_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(new_n542_), .A3(new_n779_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n781_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n782_), .A2(new_n784_), .A3(new_n547_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n767_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n758_), .B1(new_n788_), .B2(new_n629_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n777_), .A2(new_n779_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .A3(new_n778_), .A4(new_n542_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(new_n781_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n710_), .A3(new_n562_), .A4(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n766_), .B1(new_n793_), .B2(new_n786_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n786_), .A2(new_n547_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n764_), .A3(new_n780_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n796_), .A2(KEYINPUT58), .A3(new_n764_), .A4(new_n780_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n623_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n789_), .A2(new_n795_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n246_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n564_), .A2(KEYINPUT115), .A3(new_n594_), .A4(new_n245_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n710_), .B1(new_n548_), .B2(new_n563_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n806_), .B2(new_n245_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n624_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT116), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n558_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n594_), .B(new_n245_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n804_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n624_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(KEYINPUT54), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n816_), .B1(new_n815_), .B2(new_n624_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT116), .B(new_n623_), .C1(new_n814_), .C2(new_n804_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n459_), .B1(new_n803_), .B2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n316_), .A2(new_n389_), .A3(new_n634_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n710_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT121), .B1(new_n803_), .B2(new_n823_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n830_), .A2(new_n826_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n826_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n594_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n833_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g633(.A(new_n305_), .B1(new_n564_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n827_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n305_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n564_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n305_), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n827_), .B2(new_n245_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n832_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n245_), .A2(G127gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT122), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n839_), .B1(new_n840_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n827_), .B2(new_n629_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n624_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(G134gat), .ZN(G1343gat));
  AND4_X1   g645(.A1(new_n389_), .A2(new_n824_), .A3(new_n465_), .A4(new_n316_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n710_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n565_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n245_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  AOI21_X1  g653(.A(G162gat), .B1(new_n847_), .B2(new_n629_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n665_), .A2(G162gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n847_), .B2(new_n856_), .ZN(G1347gat));
  AOI21_X1  g656(.A(new_n389_), .B1(new_n803_), .B2(new_n823_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n315_), .A2(new_n459_), .A3(new_n634_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT123), .Z(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n284_), .B1(new_n862_), .B2(new_n710_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(KEYINPUT62), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n710_), .A3(new_n256_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(KEYINPUT62), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n861_), .A2(new_n564_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n257_), .ZN(G1349gat));
  NOR2_X1   g668(.A1(new_n861_), .A2(new_n246_), .ZN(new_n870_));
  MUX2_X1   g669(.A(G183gat), .B(new_n274_), .S(new_n870_), .Z(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n861_), .B2(new_n624_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n629_), .A2(new_n277_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n861_), .B2(new_n873_), .ZN(G1351gat));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n803_), .A2(new_n823_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n465_), .A2(new_n495_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n315_), .A2(new_n453_), .ZN(new_n878_));
  AND4_X1   g677(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .A4(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n803_), .B2(new_n823_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n877_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n594_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT125), .B(G197gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1352gat));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n564_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(G204gat), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(G204gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n887_), .B2(new_n889_), .ZN(G1353gat));
  OAI21_X1  g691(.A(new_n245_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n893_), .B2(new_n894_), .ZN(G1354gat));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n623_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G218gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n630_), .A2(G218gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n782_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n904_), .A2(new_n787_), .A3(new_n562_), .A4(new_n792_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n758_), .B(new_n629_), .C1(new_n905_), .C2(new_n766_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n794_), .B2(new_n630_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n245_), .B1(new_n908_), .B2(new_n801_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n818_), .A2(new_n822_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n877_), .B(new_n878_), .C1(new_n909_), .C2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT124), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n881_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n624_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n902_), .B(new_n898_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n903_), .A2(new_n917_), .ZN(G1355gat));
endmodule


