//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT36), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT68), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(KEYINPUT68), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n223_), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n212_), .A2(KEYINPUT66), .A3(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(new_n212_), .B2(new_n219_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n222_), .A2(new_n223_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT72), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G43gat), .B(G50gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  AOI21_X1  g034(.A(new_n212_), .B1(KEYINPUT9), .B2(new_n208_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n216_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(G92gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(G85gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT65), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n231_), .A2(new_n235_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n235_), .B(KEYINPUT15), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n243_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G232gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT35), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n250_), .A2(KEYINPUT35), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(KEYINPUT35), .A3(new_n250_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n207_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n256_), .A2(KEYINPUT74), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n258_), .A3(new_n255_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(KEYINPUT74), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n257_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT37), .ZN(new_n265_));
  INV_X1    g064(.A(new_n256_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n259_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT37), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G230gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  XOR2_X1   g074(.A(G71gat), .B(G78gat), .Z(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n246_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT12), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n277_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n231_), .A2(new_n243_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT12), .A3(new_n280_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n272_), .B1(new_n283_), .B2(new_n280_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT70), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G120gat), .B(G148gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G176gat), .B(G204gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n287_), .A2(new_n294_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT13), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n282_), .B(new_n300_), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT76), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(G15gat), .ZN(new_n303_));
  INV_X1    g102(.A(G22gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G1gat), .ZN(new_n306_));
  INV_X1    g105(.A(G8gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n302_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G155gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G183gat), .B(G211gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n318_), .B2(new_n312_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT78), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n298_), .A2(KEYINPUT13), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n299_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n271_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G155gat), .B(G162gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT89), .Z(new_n333_));
  OR2_X1    g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT3), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(KEYINPUT3), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(KEYINPUT2), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n337_), .B2(KEYINPUT2), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n335_), .B(new_n336_), .C1(new_n338_), .C2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT88), .Z(new_n343_));
  OAI21_X1  g142(.A(new_n333_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n334_), .A2(new_n345_), .A3(new_n339_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(KEYINPUT1), .B2(new_n332_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT28), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(KEYINPUT93), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(KEYINPUT93), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT92), .Z(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(G197gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(G197gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT21), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n362_), .B2(new_n359_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n357_), .B(new_n361_), .C1(KEYINPUT21), .C2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n356_), .B(KEYINPUT92), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n364_), .A3(KEYINPUT21), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(KEYINPUT90), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G78gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G106gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n370_), .B(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n354_), .A2(new_n355_), .A3(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n353_), .A2(KEYINPUT93), .A3(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT81), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT26), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(KEYINPUT26), .B2(new_n390_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n389_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(KEYINPUT26), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n399_), .A2(new_n396_), .A3(new_n390_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n388_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT84), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n388_), .B(new_n403_), .C1(new_n398_), .C2(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT23), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n387_), .A2(KEYINPUT24), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n406_), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT22), .ZN(new_n412_));
  OAI21_X1  g211(.A(G169gat), .B1(new_n412_), .B2(KEYINPUT85), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n385_), .A2(KEYINPUT22), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n413_), .B(new_n386_), .C1(KEYINPUT85), .C2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n415_), .A3(new_n384_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT86), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n410_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n421_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G127gat), .B(G134gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G120gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n425_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G15gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT30), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT31), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n348_), .A2(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n348_), .A2(new_n428_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT4), .A3(new_n438_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n428_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n438_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n436_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(new_n443_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G1gat), .B(G29gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT96), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT0), .B(G57gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n442_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n456_), .A2(new_n454_), .A3(new_n447_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n429_), .A2(new_n434_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n435_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT27), .ZN(new_n462_));
  INV_X1    g261(.A(new_n416_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n408_), .B1(new_n401_), .B2(KEYINPUT84), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT86), .B(new_n463_), .C1(new_n464_), .C2(new_n404_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n419_), .B1(new_n410_), .B2(new_n416_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n369_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT19), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n412_), .A2(G169gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n414_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n411_), .B(new_n384_), .C1(G176gat), .C2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(new_n387_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT26), .B(G190gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n389_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n406_), .A4(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n471_), .B1(new_n368_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n467_), .A2(new_n470_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n418_), .A2(new_n368_), .A3(new_n420_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT20), .B1(new_n368_), .B2(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n470_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G8gat), .B(G36gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n483_), .A2(new_n487_), .A3(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n465_), .A2(new_n466_), .A3(new_n369_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n469_), .B1(new_n495_), .B2(new_n485_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n467_), .A2(new_n470_), .A3(new_n482_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n462_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT100), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n492_), .A3(new_n497_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT100), .A3(new_n462_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n495_), .A2(new_n469_), .A3(new_n485_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n470_), .B1(new_n467_), .B2(new_n482_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n493_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n509_), .A2(KEYINPUT27), .A3(new_n503_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT101), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT101), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n513_), .B(new_n510_), .C1(new_n501_), .C2(new_n505_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n381_), .B(new_n461_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT102), .ZN(new_n516_));
  INV_X1    g315(.A(new_n381_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT100), .B1(new_n504_), .B2(new_n462_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n500_), .B(KEYINPUT27), .C1(new_n502_), .C2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n513_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n511_), .B(KEYINPUT101), .C1(new_n518_), .C2(new_n519_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT102), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n461_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n492_), .A2(KEYINPUT32), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT98), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n496_), .A2(new_n497_), .A3(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n458_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT99), .ZN(new_n531_));
  OR2_X1    g330(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n454_), .B(new_n532_), .C1(new_n456_), .C2(new_n447_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n454_), .B1(new_n446_), .B2(new_n443_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  OR3_X1    g336(.A1(new_n533_), .A2(new_n537_), .A3(new_n504_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n458_), .A2(new_n539_), .A3(new_n529_), .A4(new_n528_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n381_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n517_), .A2(new_n459_), .A3(new_n506_), .A4(new_n511_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n435_), .A2(new_n460_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n516_), .A2(new_n525_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n311_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n245_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n311_), .B2(new_n235_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n311_), .B(new_n235_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n548_), .A2(new_n551_), .B1(new_n552_), .B2(new_n550_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT80), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n553_), .A2(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n546_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n331_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT103), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT103), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n331_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n459_), .A2(G1gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n202_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n202_), .A3(new_n568_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT38), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n567_), .A2(new_n202_), .A3(new_n568_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n544_), .A2(new_n545_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n521_), .A2(new_n522_), .ZN(new_n577_));
  AND4_X1   g376(.A1(new_n524_), .A2(new_n577_), .A3(new_n381_), .A4(new_n461_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n524_), .B1(new_n523_), .B2(new_n461_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n267_), .A2(KEYINPUT105), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n267_), .A2(KEYINPUT105), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n580_), .A2(KEYINPUT106), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT106), .B1(new_n580_), .B2(new_n584_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n299_), .A2(new_n327_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(new_n561_), .A3(new_n325_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n458_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(G1gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n572_), .A2(new_n575_), .A3(new_n592_), .ZN(G1324gat));
  INV_X1    g392(.A(new_n577_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n567_), .A2(new_n307_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n594_), .B(new_n590_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(G8gat), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n597_), .A2(new_n596_), .A3(G8gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n595_), .B(KEYINPUT40), .C1(new_n598_), .C2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1325gat));
  INV_X1    g403(.A(new_n545_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n567_), .A2(new_n431_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n587_), .A2(new_n605_), .A3(new_n590_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n607_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(new_n607_), .B2(G15gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(G1326gat));
  NAND3_X1  g409(.A1(new_n567_), .A2(new_n304_), .A3(new_n517_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n587_), .A2(new_n517_), .A3(new_n590_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G22gat), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(G1327gat));
  NAND2_X1  g415(.A1(new_n583_), .A2(new_n325_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT109), .Z(new_n618_));
  AND3_X1   g417(.A1(new_n562_), .A2(new_n588_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G29gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n458_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT107), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n265_), .A2(new_n622_), .A3(new_n269_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT43), .B1(new_n546_), .B2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n270_), .A2(KEYINPUT43), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n580_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n588_), .A2(new_n560_), .A3(new_n325_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT44), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n634_), .B(new_n631_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n458_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n637_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT108), .B1(new_n637_), .B2(G29gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n621_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n619_), .A2(new_n641_), .A3(new_n594_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n633_), .A2(new_n635_), .A3(new_n577_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT46), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n643_), .B(KEYINPUT46), .C1(new_n641_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1329gat));
  AOI21_X1  g448(.A(G43gat), .B1(new_n619_), .B2(new_n605_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n545_), .A2(new_n423_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n636_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g452(.A(G50gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n619_), .A2(new_n654_), .A3(new_n517_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT110), .B1(new_n636_), .B2(new_n517_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n625_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n623_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n580_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n628_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n546_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n632_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n634_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n632_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(KEYINPUT110), .A3(new_n517_), .A4(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G50gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n655_), .B1(new_n656_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT111), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT111), .B(new_n655_), .C1(new_n656_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1331gat));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n546_), .A2(new_n560_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n271_), .A2(new_n325_), .A3(new_n588_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(new_n459_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT112), .Z(new_n678_));
  AND4_X1   g477(.A1(new_n561_), .A2(new_n587_), .A3(new_n326_), .A4(new_n589_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n459_), .A2(new_n673_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(G1332gat));
  INV_X1    g480(.A(new_n676_), .ZN(new_n682_));
  INV_X1    g481(.A(G64gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n594_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n594_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G64gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT48), .B(new_n683_), .C1(new_n679_), .C2(new_n594_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(KEYINPUT49), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n679_), .A2(new_n605_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(G71gat), .ZN(new_n692_));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT49), .B(new_n693_), .C1(new_n679_), .C2(new_n605_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n605_), .A2(new_n693_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT113), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n692_), .A2(new_n694_), .B1(new_n676_), .B2(new_n696_), .ZN(G1334gat));
  INV_X1    g496(.A(G78gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n682_), .A2(new_n698_), .A3(new_n517_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT50), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n679_), .A2(new_n517_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(G78gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT50), .B(new_n698_), .C1(new_n679_), .C2(new_n517_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1335gat));
  AND3_X1   g503(.A1(new_n674_), .A2(new_n589_), .A3(new_n618_), .ZN(new_n705_));
  INV_X1    g504(.A(G85gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n458_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n588_), .A2(new_n560_), .A3(new_n326_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n630_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT114), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n458_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n712_), .B2(new_n706_), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n705_), .B2(new_n594_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n594_), .A2(new_n239_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n711_), .B2(new_n715_), .ZN(G1337gat));
  AOI21_X1  g515(.A(new_n215_), .B1(new_n709_), .B2(new_n605_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n705_), .A2(new_n605_), .A3(new_n237_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n718_), .B1(new_n719_), .B2(KEYINPUT51), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT51), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n705_), .A2(new_n216_), .A3(new_n517_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT116), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n630_), .A2(new_n517_), .A3(new_n708_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .A4(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n216_), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n725_), .A2(new_n728_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n723_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT54), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n329_), .B2(new_n561_), .ZN(new_n733_));
  NOR4_X1   g532(.A1(new_n271_), .A2(new_n328_), .A3(KEYINPUT54), .A4(new_n560_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n560_), .A2(new_n295_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n285_), .B(KEYINPUT55), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n281_), .A2(new_n273_), .A3(new_n284_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT117), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n281_), .A2(new_n284_), .A3(new_n740_), .A4(new_n273_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n294_), .B1(new_n737_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n285_), .A2(KEYINPUT55), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n285_), .A2(KEYINPUT55), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n293_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT119), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n744_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n747_), .A2(new_n293_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n747_), .C2(new_n293_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n736_), .B1(new_n751_), .B2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n552_), .A2(new_n549_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n759_), .A2(new_n556_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT120), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n549_), .B1(new_n311_), .B2(new_n235_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n760_), .A2(new_n761_), .B1(new_n548_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n761_), .B2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n558_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n298_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT57), .B(new_n584_), .C1(new_n758_), .C2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT118), .B1(new_n743_), .B2(KEYINPUT56), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n753_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n744_), .A3(new_n770_), .A4(new_n750_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n736_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n766_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(new_n583_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n765_), .A2(new_n296_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n753_), .A2(new_n754_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n748_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n271_), .B1(new_n778_), .B2(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n748_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n775_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT121), .B1(new_n779_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n782_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(KEYINPUT58), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .A4(new_n271_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n767_), .A2(new_n774_), .A3(new_n784_), .A4(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n735_), .B1(new_n789_), .B2(new_n325_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n523_), .A2(new_n458_), .A3(new_n605_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n560_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n271_), .A3(new_n787_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n767_), .A2(new_n774_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n325_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n735_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n792_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n796_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n561_), .A2(KEYINPUT122), .ZN(new_n805_));
  MUX2_X1   g604(.A(KEYINPUT122), .B(new_n805_), .S(G113gat), .Z(new_n806_));
  AOI21_X1  g605(.A(new_n795_), .B1(new_n804_), .B2(new_n806_), .ZN(G1340gat));
  NAND3_X1  g606(.A1(new_n796_), .A2(new_n589_), .A3(new_n803_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G120gat), .ZN(new_n809_));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n794_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1341gat));
  NAND3_X1  g612(.A1(new_n796_), .A2(new_n326_), .A3(new_n803_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G127gat), .ZN(new_n815_));
  OR3_X1    g614(.A1(new_n793_), .A2(G127gat), .A3(new_n325_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1342gat));
  NAND3_X1  g616(.A1(new_n796_), .A2(new_n271_), .A3(new_n803_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G134gat), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n793_), .A2(G134gat), .A3(new_n584_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1343gat));
  NOR2_X1   g620(.A1(new_n790_), .A2(new_n605_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n594_), .A2(new_n459_), .A3(new_n381_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n560_), .A3(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT123), .B(G141gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1344gat));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n589_), .A3(new_n823_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n326_), .A3(new_n823_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AND2_X1   g630(.A1(new_n822_), .A2(new_n823_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G162gat), .B1(new_n832_), .B2(new_n583_), .ZN(new_n833_));
  INV_X1    g632(.A(G162gat), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n626_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n832_), .B2(new_n835_), .ZN(G1347gat));
  AOI21_X1  g635(.A(new_n735_), .B1(new_n798_), .B2(new_n325_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n517_), .A2(new_n545_), .A3(new_n458_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n594_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n560_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n385_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n841_), .B(new_n842_), .C1(KEYINPUT124), .C2(KEYINPUT62), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n845_), .B(new_n846_), .C1(new_n473_), .C2(new_n841_), .ZN(G1348gat));
  NOR2_X1   g646(.A1(new_n588_), .A2(new_n386_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n790_), .A2(new_n839_), .A3(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n837_), .A2(new_n588_), .A3(new_n839_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n850_), .A2(KEYINPUT125), .B1(new_n851_), .B2(G176gat), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n850_), .A2(KEYINPUT125), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT126), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n850_), .A2(KEYINPUT125), .ZN(new_n855_));
  INV_X1    g654(.A(new_n839_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n801_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n386_), .B1(new_n857_), .B2(new_n588_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(KEYINPUT125), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n855_), .A2(new_n858_), .A3(new_n859_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n854_), .A2(new_n861_), .ZN(G1349gat));
  NOR3_X1   g661(.A1(new_n857_), .A2(new_n389_), .A3(new_n325_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n790_), .A2(new_n839_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G183gat), .B1(new_n864_), .B2(new_n326_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n857_), .B2(new_n270_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n840_), .A2(new_n478_), .A3(new_n583_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1351gat));
  NOR3_X1   g668(.A1(new_n577_), .A2(new_n458_), .A3(new_n381_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n822_), .A2(new_n560_), .A3(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g671(.A1(new_n822_), .A2(new_n870_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n588_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT127), .B(G204gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1353gat));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n325_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT63), .B(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n877_), .B2(new_n880_), .ZN(G1354gat));
  OAI21_X1  g680(.A(G218gat), .B1(new_n873_), .B2(new_n270_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n584_), .A2(G218gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n873_), .B2(new_n883_), .ZN(G1355gat));
endmodule


