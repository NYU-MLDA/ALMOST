//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT74), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n211_), .B(KEYINPUT14), .C1(new_n207_), .C2(new_n208_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n206_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G229gat), .A2(G233gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n206_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n216_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(new_n216_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n219_), .B1(new_n223_), .B2(new_n218_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G197gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n218_), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n232_), .B(new_n221_), .C1(new_n222_), .C2(new_n216_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n233_), .B2(new_n219_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT76), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n228_), .ZN(new_n238_));
  INV_X1    g037(.A(G204gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT82), .A2(G197gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n228_), .A2(G204gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n238_), .A2(KEYINPUT83), .A3(new_n239_), .A4(new_n240_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT21), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n228_), .A2(G204gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n238_), .A2(new_n240_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT21), .B(new_n249_), .C1(new_n250_), .C2(G204gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT25), .B(G183gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n255_));
  INV_X1    g054(.A(G190gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(KEYINPUT26), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G190gat), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n254_), .B(new_n257_), .C1(new_n258_), .C2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n226_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT24), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n226_), .A3(new_n265_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n259_), .A2(new_n264_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n265_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT78), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT22), .B(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n265_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n262_), .B(new_n263_), .C1(G183gat), .C2(G190gat), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n267_), .A4(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n271_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n249_), .B1(new_n250_), .B2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n248_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(KEYINPUT21), .C1(new_n283_), .C2(new_n282_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n253_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n251_), .B1(new_n246_), .B2(KEYINPUT21), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  INV_X1    g087(.A(new_n282_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(KEYINPUT84), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n287_), .A2(new_n248_), .B1(new_n290_), .B2(new_n284_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n269_), .A2(KEYINPUT87), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT24), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n294_), .A3(new_n267_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(KEYINPUT88), .A3(new_n267_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(new_n266_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n264_), .B(new_n301_), .C1(new_n266_), .C2(new_n298_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n266_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n262_), .A2(new_n263_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT89), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n254_), .A2(new_n258_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n279_), .A2(new_n267_), .A3(new_n274_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n286_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n253_), .A2(new_n285_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n271_), .A2(new_n280_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n291_), .A2(new_n309_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(KEYINPUT90), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n317_), .A2(new_n322_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT18), .B(G64gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G92gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n323_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(KEYINPUT91), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n324_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n338_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(KEYINPUT2), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(KEYINPUT81), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n337_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n353_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  OAI221_X1 g153(.A(new_n354_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n336_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT79), .B(G127gat), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G134gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(G113gat), .B(G120gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(G127gat), .ZN(new_n359_));
  INV_X1    g158(.A(G134gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n360_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n352_), .A2(new_n355_), .A3(new_n362_), .A4(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n362_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n339_), .A2(new_n340_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n369_), .A2(new_n351_), .A3(new_n344_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n355_), .B1(new_n370_), .B2(new_n336_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n372_), .A3(KEYINPUT92), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT4), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT93), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n372_), .A2(KEYINPUT4), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n378_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G1gat), .B(G29gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT95), .ZN(new_n385_));
  XOR2_X1   g184(.A(G57gat), .B(G85gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND3_X1  g188(.A1(new_n382_), .A2(new_n383_), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n376_), .A2(new_n380_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n382_), .A2(KEYINPUT33), .A3(new_n383_), .A4(new_n389_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT96), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n335_), .A2(new_n392_), .A3(new_n396_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n328_), .A2(KEYINPUT32), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT98), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n324_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n310_), .A2(new_n312_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n318_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n390_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n389_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n408_));
  OAI221_X1 g207(.A(new_n403_), .B1(new_n406_), .B2(new_n401_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n316_), .B(KEYINPUT30), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n368_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT30), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n281_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n316_), .A2(KEYINPUT30), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n418_), .A2(new_n362_), .A3(new_n366_), .A4(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n414_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n416_), .A2(new_n420_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n422_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n413_), .A3(new_n424_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n427_), .A2(new_n430_), .A3(KEYINPUT80), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT80), .B1(new_n427_), .B2(new_n430_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n315_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n315_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n434_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(G50gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(G50gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT28), .B(G22gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n452_), .A3(new_n448_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n442_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n439_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n437_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT86), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n445_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n451_), .A2(new_n453_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n434_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n410_), .A2(new_n433_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n332_), .A2(new_n465_), .A3(new_n334_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT100), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n332_), .A2(KEYINPUT100), .A3(new_n465_), .A4(new_n334_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n329_), .B(KEYINPUT27), .C1(new_n328_), .C2(new_n406_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n408_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT99), .A3(new_n390_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n460_), .B(new_n462_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n427_), .A2(new_n430_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n463_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n470_), .A2(new_n471_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n236_), .B1(new_n464_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT7), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT6), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  AOI21_X1  g288(.A(new_n483_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT66), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n487_), .B(KEYINPUT65), .ZN(new_n492_));
  INV_X1    g291(.A(new_n485_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n483_), .B(new_n489_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(KEYINPUT66), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n491_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G85gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(G85gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(G92gat), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT10), .B(G99gat), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n501_), .B(new_n502_), .C1(G106gat), .C2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n492_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n222_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n490_), .B(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n510_), .B2(new_n494_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n206_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n516_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n515_), .A2(new_n516_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n508_), .A2(new_n512_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT72), .B(G134gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G162gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G190gat), .B(G218gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT36), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n517_), .A2(new_n520_), .A3(KEYINPUT73), .A4(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n517_), .A2(new_n520_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n524_), .B(KEYINPUT36), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n531_), .A2(KEYINPUT37), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT37), .B1(new_n531_), .B2(new_n534_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n542_), .A3(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n216_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549_));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n548_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(KEYINPUT17), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n538_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT67), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n511_), .B2(new_n545_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n545_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n507_), .A2(new_n564_), .B1(KEYINPUT67), .B2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(KEYINPUT67), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n545_), .B(new_n566_), .C1(new_n496_), .C2(new_n506_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n562_), .B(new_n563_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n511_), .A2(new_n545_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n507_), .A2(new_n564_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n239_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n265_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT13), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT68), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n482_), .A2(new_n559_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n207_), .A3(new_n476_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT101), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n531_), .A2(new_n534_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n591_), .B(new_n558_), .C1(new_n464_), .C2(new_n481_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n582_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n235_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n476_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n589_), .A3(new_n599_), .ZN(G1324gat));
  NAND2_X1  g399(.A1(new_n470_), .A2(new_n471_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n584_), .A2(new_n208_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n601_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(G8gat), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT39), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT39), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n597_), .B2(new_n433_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT102), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT41), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n610_), .B(KEYINPUT102), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT41), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n433_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n584_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n615_), .A3(new_n618_), .ZN(G1326gat));
  INV_X1    g418(.A(G22gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n463_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n596_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n584_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  NOR2_X1   g424(.A1(new_n590_), .A2(new_n557_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n482_), .A2(new_n582_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n476_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n593_), .A2(new_n594_), .A3(new_n557_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n464_), .A2(new_n481_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(new_n538_), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT43), .B(new_n537_), .C1(new_n464_), .C2(new_n481_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT44), .B(new_n629_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(new_n476_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n628_), .B1(new_n639_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n627_), .A2(new_n641_), .A3(new_n601_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n601_), .A3(new_n637_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n644_), .B2(G36gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n643_), .B(KEYINPUT46), .C1(new_n645_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  NAND3_X1  g450(.A1(new_n638_), .A2(G43gat), .A3(new_n478_), .ZN(new_n652_));
  INV_X1    g451(.A(G43gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n627_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n433_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g456(.A(G50gat), .B1(new_n627_), .B2(new_n621_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n621_), .A2(G50gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n638_), .B2(new_n659_), .ZN(G1331gat));
  AOI21_X1  g459(.A(new_n235_), .B1(new_n464_), .B2(new_n481_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(new_n593_), .A3(new_n559_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G57gat), .B1(new_n662_), .B2(new_n476_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n583_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n592_), .A2(new_n236_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(G57gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(KEYINPUT104), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  OAI21_X1  g468(.A(G57gat), .B1(new_n598_), .B2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n663_), .B1(new_n668_), .B2(new_n670_), .ZN(G1332gat));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n665_), .B2(new_n601_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n662_), .A2(new_n672_), .A3(new_n601_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n665_), .B2(new_n617_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT49), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n662_), .A2(new_n677_), .A3(new_n617_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1334gat));
  INV_X1    g480(.A(G78gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n662_), .A2(new_n682_), .A3(new_n621_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G78gat), .B1(new_n666_), .B2(new_n463_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT50), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT50), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT105), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n683_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1335gat));
  NAND3_X1  g490(.A1(new_n664_), .A2(new_n626_), .A3(new_n661_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n476_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n632_), .A2(new_n633_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n557_), .A2(new_n235_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n593_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n500_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n598_), .B2(new_n498_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n694_), .B1(new_n701_), .B2(new_n703_), .ZN(G1336gat));
  NAND2_X1  g503(.A1(new_n601_), .A2(G92gat), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT107), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n601_), .ZN(new_n709_));
  INV_X1    g508(.A(G92gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n708_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n706_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n697_), .B2(new_n433_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n503_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n693_), .A2(new_n478_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g521(.A1(new_n695_), .A2(new_n621_), .A3(new_n593_), .A4(new_n696_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(G106gat), .A3(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n692_), .A2(G106gat), .A3(new_n463_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n723_), .A2(G106gat), .A3(new_n729_), .A4(new_n724_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n727_), .A2(new_n733_), .A3(new_n728_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1339gat));
  XOR2_X1   g534(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n568_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n566_), .B1(new_n511_), .B2(new_n545_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n507_), .A2(KEYINPUT67), .A3(new_n560_), .A4(new_n564_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT112), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n740_), .A2(new_n563_), .A3(new_n562_), .A4(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n562_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n569_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n737_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n578_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n578_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(KEYINPUT113), .A3(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n750_), .A2(KEYINPUT113), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n235_), .A2(KEYINPUT111), .A3(new_n580_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT111), .B1(new_n235_), .B2(new_n580_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n217_), .A2(new_n232_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n223_), .B(KEYINPUT114), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n229_), .B(new_n757_), .C1(new_n758_), .C2(new_n218_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n231_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n581_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT57), .A3(new_n590_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n750_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n578_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n580_), .B(new_n760_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n749_), .A2(new_n750_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n580_), .A4(new_n760_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n538_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n591_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n763_), .B(new_n771_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n558_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n536_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n531_), .A2(KEYINPUT37), .A3(new_n534_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n594_), .A2(KEYINPUT76), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT76), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n235_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n778_), .A2(KEYINPUT110), .A3(new_n780_), .A4(new_n557_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n776_), .A2(new_n777_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT110), .B1(new_n236_), .B2(new_n557_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n582_), .A4(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n776_), .A2(new_n582_), .A3(new_n777_), .A4(new_n781_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT54), .B1(new_n787_), .B2(new_n784_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n601_), .A2(new_n598_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n479_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(KEYINPUT117), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n789_), .B1(new_n774_), .B2(new_n558_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n797_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n235_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n797_), .A2(KEYINPUT59), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .B1(KEYINPUT57), .B2(new_n772_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n771_), .B(new_n808_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n557_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n810_), .B2(new_n789_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT59), .B1(new_n801_), .B2(new_n797_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n236_), .A2(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT119), .Z(new_n816_));
  AOI21_X1  g615(.A(new_n804_), .B1(new_n813_), .B2(new_n816_), .ZN(G1340gat));
  NAND2_X1  g616(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n763_), .A3(new_n809_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n789_), .B1(new_n819_), .B2(new_n558_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n797_), .A2(KEYINPUT59), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n812_), .B(new_n664_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n811_), .A2(KEYINPUT120), .A3(new_n664_), .A4(new_n812_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(G120gat), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n803_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(G1341gat));
  XNOR2_X1  g629(.A(KEYINPUT122), .B(G127gat), .ZN(new_n831_));
  AND4_X1   g630(.A1(new_n557_), .A2(new_n811_), .A3(new_n812_), .A4(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n803_), .A2(new_n557_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n558_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT121), .B1(new_n837_), .B2(G127gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n836_), .B2(new_n838_), .ZN(G1342gat));
  AOI21_X1  g638(.A(G134gat), .B1(new_n803_), .B2(new_n591_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n538_), .A2(G134gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT123), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n813_), .B2(new_n842_), .ZN(G1343gat));
  NOR4_X1   g642(.A1(new_n801_), .A2(new_n601_), .A3(new_n598_), .A4(new_n477_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n235_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n664_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n557_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT124), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n849_), .B(new_n851_), .ZN(G1346gat));
  INV_X1    g651(.A(G162gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n844_), .B2(new_n538_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n801_), .A2(new_n477_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n590_), .A2(G162gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n855_), .A2(new_n792_), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT125), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n792_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G162gat), .B1(new_n859_), .B2(new_n537_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n844_), .A2(new_n856_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(G1347gat));
  AOI21_X1  g663(.A(new_n476_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(new_n617_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n463_), .B(new_n866_), .C1(new_n810_), .C2(new_n789_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G169gat), .B1(new_n867_), .B2(new_n594_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n867_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n235_), .A3(new_n276_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT62), .B(G169gat), .C1(new_n867_), .C2(new_n594_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(G1348gat));
  AOI21_X1  g673(.A(G176gat), .B1(new_n871_), .B2(new_n593_), .ZN(new_n875_));
  OR3_X1    g674(.A1(new_n801_), .A2(KEYINPUT126), .A3(new_n621_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT126), .B1(new_n801_), .B2(new_n621_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n265_), .B(new_n583_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n866_), .B2(new_n878_), .ZN(G1349gat));
  NOR3_X1   g678(.A1(new_n867_), .A2(new_n254_), .A3(new_n558_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n877_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n557_), .A3(new_n866_), .ZN(new_n882_));
  INV_X1    g681(.A(G183gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n882_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n867_), .B2(new_n537_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n591_), .A2(new_n258_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n867_), .B2(new_n886_), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n855_), .A2(new_n865_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n594_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n228_), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n583_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n239_), .ZN(G1353gat));
  NAND3_X1  g691(.A1(new_n855_), .A2(new_n557_), .A3(new_n865_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n893_), .B2(new_n894_), .ZN(G1354gat));
  NOR2_X1   g696(.A1(new_n888_), .A2(new_n590_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G218gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n888_), .A2(new_n537_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(G218gat), .B2(new_n900_), .ZN(G1355gat));
endmodule


