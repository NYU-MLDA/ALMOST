//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G120gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G113gat), .ZN(new_n209_));
  INV_X1    g008(.A(G113gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G120gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n207_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(new_n212_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT88), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n207_), .A2(new_n212_), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n204_), .A2(new_n206_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT31), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(new_n223_), .B2(KEYINPUT82), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(G190gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(KEYINPUT24), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n228_), .A2(new_n233_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G169gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n231_), .B(new_n232_), .C1(G183gat), .C2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT83), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT30), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(G71gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G99gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G15gat), .B(G43gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT87), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n259_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n240_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n247_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT30), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n202_), .B(new_n221_), .C1(new_n262_), .C2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n268_), .B(KEYINPUT86), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n261_), .B(KEYINPUT87), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n221_), .A2(new_n202_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n221_), .A2(new_n202_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G85gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n283_));
  OR2_X1    g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT90), .B1(new_n282_), .B2(KEYINPUT1), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT91), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(KEYINPUT1), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(KEYINPUT1), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n284_), .A4(new_n283_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n217_), .A2(new_n218_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n284_), .A2(new_n282_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n298_), .B(KEYINPUT3), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n296_), .B(KEYINPUT2), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n215_), .A2(new_n219_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n306_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n309_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT101), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n299_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n285_), .A2(new_n286_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n288_), .B1(new_n316_), .B2(new_n293_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n317_), .B2(new_n287_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n220_), .B1(new_n318_), .B2(new_n306_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT101), .A3(new_n309_), .A4(new_n308_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n311_), .A2(new_n310_), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n306_), .B(new_n301_), .C1(new_n295_), .C2(new_n299_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT4), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n309_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n281_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n309_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n325_), .B1(new_n319_), .B2(new_n308_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n322_), .A2(KEYINPUT4), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n281_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n314_), .A4(new_n320_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n277_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n300_), .A2(new_n307_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT96), .ZN(new_n339_));
  INV_X1    g138(.A(G218gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G211gat), .ZN(new_n341_));
  INV_X1    g140(.A(G211gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G218gat), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n341_), .A2(new_n343_), .A3(KEYINPUT95), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT95), .B1(new_n341_), .B2(new_n343_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n339_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT94), .B(G204gat), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n347_), .B(new_n348_), .C1(new_n349_), .C2(G197gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT95), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n342_), .A2(G218gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n340_), .A2(G211gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n341_), .A2(new_n343_), .A3(KEYINPUT95), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT96), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n346_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n355_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n347_), .B1(G197gat), .B2(G204gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n349_), .B2(G197gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n348_), .B1(new_n349_), .B2(G197gat), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n358_), .B(new_n360_), .C1(KEYINPUT21), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT97), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT97), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT93), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n338_), .A2(new_n363_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n367_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n338_), .A2(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n372_), .A2(KEYINPUT98), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT98), .B1(new_n372_), .B2(new_n374_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n311_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(KEYINPUT28), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(KEYINPUT28), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(new_n374_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n375_), .A2(new_n376_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT92), .B1(new_n384_), .B2(new_n385_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n385_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n383_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n372_), .A2(new_n374_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n389_), .B(new_n392_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT106), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n236_), .A2(new_n237_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT100), .B(KEYINPUT24), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT26), .B(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n222_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n400_), .A2(new_n233_), .A3(new_n401_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n244_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n363_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT20), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT105), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n364_), .A2(new_n249_), .A3(new_n366_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(KEYINPUT105), .A3(KEYINPUT20), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT19), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n249_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT99), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n363_), .A2(new_n405_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n357_), .A2(new_n365_), .A3(new_n362_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n365_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n266_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT99), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT20), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n415_), .B1(new_n414_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT18), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n424_), .A2(new_n419_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n423_), .B1(new_n422_), .B2(KEYINPUT20), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n414_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n414_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n436_), .A4(new_n406_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n430_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(KEYINPUT27), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT27), .ZN(new_n440_));
  INV_X1    g239(.A(new_n437_), .ZN(new_n441_));
  AOI211_X1 g240(.A(new_n431_), .B(new_n441_), .C1(new_n425_), .C2(new_n414_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n430_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n440_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n397_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n439_), .A2(new_n397_), .A3(new_n444_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n336_), .B(new_n396_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n335_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n448_), .A2(new_n444_), .A3(new_n439_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT103), .ZN(new_n450_));
  INV_X1    g249(.A(new_n419_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n364_), .A2(new_n366_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n417_), .B1(new_n452_), .B2(new_n266_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n453_), .B2(new_n423_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n436_), .B1(new_n454_), .B2(new_n418_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n431_), .B1(new_n455_), .B2(new_n441_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n329_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n322_), .A2(new_n323_), .A3(new_n309_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n457_), .A2(new_n333_), .A3(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n321_), .A2(new_n327_), .A3(new_n281_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(KEYINPUT33), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n461_), .A3(new_n438_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n334_), .A2(KEYINPUT102), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT102), .B1(new_n334_), .B2(new_n463_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n450_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n442_), .A2(new_n443_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n460_), .B2(KEYINPUT33), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n334_), .A2(KEYINPUT102), .A3(new_n463_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n468_), .A2(new_n472_), .A3(KEYINPUT103), .A4(new_n461_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n426_), .A2(KEYINPUT32), .A3(new_n430_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT104), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n435_), .A2(new_n437_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(new_n335_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n467_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n449_), .B1(new_n479_), .B2(new_n396_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n277_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n447_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483_));
  INV_X1    g282(.A(G1gat), .ZN(new_n484_));
  INV_X1    g283(.A(G8gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT14), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G8gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n489_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n492_), .B(KEYINPUT15), .ZN(new_n496_));
  INV_X1    g295(.A(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n493_), .A2(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT80), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT81), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n482_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G230gat), .ZN(new_n508_));
  INV_X1    g307(.A(G233gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT10), .B(G99gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT64), .ZN(new_n513_));
  OR2_X1    g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n515_));
  NAND2_X1  g314(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT6), .ZN(new_n522_));
  INV_X1    g321(.A(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(G92gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(KEYINPUT9), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT65), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT9), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n527_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n520_), .B(new_n522_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n525_), .A2(new_n526_), .ZN(new_n533_));
  OR3_X1    g332(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT8), .B(new_n533_), .C1(new_n535_), .C2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n533_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n532_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT67), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n532_), .A2(new_n542_), .A3(new_n545_), .A4(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT11), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT69), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n548_), .B(KEYINPUT68), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n511_), .B1(new_n547_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n560_), .A2(new_n561_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(KEYINPUT70), .A3(new_n544_), .A4(new_n546_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n547_), .A2(new_n562_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n564_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n510_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n544_), .A2(new_n546_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n572_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n547_), .A2(new_n562_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n571_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n544_), .A2(new_n492_), .A3(new_n546_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT74), .A3(KEYINPUT35), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(KEYINPUT35), .B2(new_n595_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n543_), .B2(new_n496_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT74), .B1(new_n595_), .B2(KEYINPUT35), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n608_));
  OR4_X1    g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n607_), .A4(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n611_), .B2(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n609_), .A2(KEYINPUT76), .A3(new_n618_), .A4(new_n610_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n614_), .A2(new_n615_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT78), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT17), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n562_), .B(new_n489_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT77), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n629_), .B(new_n631_), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n628_), .B(new_n632_), .C1(new_n627_), .C2(new_n625_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n620_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n507_), .A2(new_n591_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n484_), .A3(new_n335_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n611_), .B(KEYINPUT107), .Z(new_n642_));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n482_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n591_), .A2(new_n506_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(new_n635_), .A3(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n335_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n640_), .B(new_n641_), .C1(new_n484_), .C2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1324gat));
  NOR2_X1   g450(.A1(new_n446_), .A2(new_n445_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n637_), .A2(new_n485_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n647_), .A2(new_n652_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(G8gat), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT39), .B(new_n485_), .C1(new_n647_), .C2(new_n652_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n658_), .B(new_n659_), .Z(G1325gat));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n647_), .B2(new_n481_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT41), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n637_), .A2(new_n661_), .A3(new_n481_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n396_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n647_), .B2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n666_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT111), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n637_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(G1327gat));
  OR2_X1    g472(.A1(new_n642_), .A2(new_n634_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n590_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n507_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n335_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n482_), .A2(new_n620_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n482_), .A2(new_n681_), .A3(new_n620_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n646_), .A2(new_n634_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n335_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n678_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n687_), .A2(new_n652_), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n652_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n676_), .A2(G36gat), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(KEYINPUT46), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  NAND4_X1  g501(.A1(new_n687_), .A2(G43gat), .A3(new_n481_), .A4(new_n688_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n676_), .A2(new_n277_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(G43gat), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g505(.A1(new_n676_), .A2(G50gat), .A3(new_n396_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n687_), .A2(new_n667_), .A3(new_n688_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT113), .ZN(new_n709_));
  OAI21_X1  g508(.A(G50gat), .B1(new_n708_), .B2(KEYINPUT113), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(G1331gat));
  INV_X1    g510(.A(new_n506_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n482_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n590_), .A3(new_n636_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT114), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n335_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(KEYINPUT115), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT115), .B1(new_n716_), .B2(new_n717_), .ZN(new_n719_));
  NOR4_X1   g518(.A1(new_n645_), .A2(new_n506_), .A3(new_n591_), .A4(new_n635_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(G57gat), .A3(new_n335_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT116), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n718_), .A2(new_n719_), .A3(new_n722_), .ZN(G1332gat));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n720_), .B2(new_n652_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT48), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n715_), .A2(new_n724_), .A3(new_n652_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1333gat));
  AOI21_X1  g527(.A(new_n252_), .B1(new_n720_), .B2(new_n481_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n715_), .A2(new_n252_), .A3(new_n481_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n720_), .B2(new_n667_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT50), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n715_), .A2(new_n733_), .A3(new_n667_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n591_), .A2(new_n506_), .A3(new_n634_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n335_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n482_), .A2(new_n712_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n591_), .A3(new_n674_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n523_), .A3(new_n335_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1336gat));
  OAI21_X1  g549(.A(G92gat), .B1(new_n744_), .B2(new_n694_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n748_), .A2(new_n524_), .A3(new_n652_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1337gat));
  OR2_X1    g552(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n754_));
  OAI21_X1  g553(.A(G99gat), .B1(new_n744_), .B2(new_n277_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n277_), .B1(new_n517_), .B2(new_n513_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n748_), .A2(new_n756_), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n277_), .B1(new_n759_), .B2(new_n741_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n754_), .B(new_n757_), .C1(new_n760_), .C2(new_n254_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n758_), .A2(new_n762_), .ZN(G1338gat));
  AND3_X1   g562(.A1(new_n482_), .A2(new_n681_), .A3(new_n620_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n681_), .B1(new_n482_), .B2(new_n620_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n667_), .B(new_n738_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G106gat), .B1(new_n766_), .B2(KEYINPUT119), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n740_), .B2(new_n667_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n740_), .A2(new_n768_), .A3(new_n667_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(KEYINPUT119), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .A4(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n748_), .A2(new_n519_), .A3(new_n667_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT124), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n636_), .A2(new_n712_), .A3(new_n591_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n500_), .A2(new_n504_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n504_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n494_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n498_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT120), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n791_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n571_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n563_), .A2(new_n566_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n510_), .B1(new_n797_), .B2(new_n576_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n577_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n568_), .A2(new_n574_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT55), .A4(new_n572_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n583_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n583_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n506_), .B(new_n796_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n793_), .A2(new_n795_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n642_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n796_), .A2(new_n791_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n814_), .A2(new_n815_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT121), .B1(new_n796_), .B2(new_n791_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT122), .A3(new_n620_), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n816_), .A2(new_n813_), .A3(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT122), .B1(new_n818_), .B2(new_n620_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n811_), .B(new_n812_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n634_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n818_), .A2(new_n620_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n820_), .A3(new_n819_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT123), .A3(new_n811_), .A4(new_n812_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n785_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n652_), .A2(new_n667_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n335_), .A3(new_n481_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n831_), .A2(new_n712_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n782_), .B1(new_n834_), .B2(G113gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n823_), .A2(new_n824_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n837_), .A2(new_n635_), .A3(new_n830_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n785_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT124), .B(new_n210_), .C1(new_n839_), .C2(new_n712_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n823_), .A2(new_n635_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n836_), .C1(new_n842_), .C2(new_n785_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n839_), .B2(KEYINPUT59), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n712_), .A2(new_n210_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n835_), .A2(new_n840_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n831_), .A2(new_n833_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n590_), .B(new_n843_), .C1(new_n848_), .C2(new_n841_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n208_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n848_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n208_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1341gat));
  OAI211_X1 g652(.A(new_n634_), .B(new_n843_), .C1(new_n848_), .C2(new_n841_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n848_), .A2(new_n205_), .A3(new_n634_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1342gat));
  OAI211_X1 g656(.A(new_n620_), .B(new_n843_), .C1(new_n848_), .C2(new_n841_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G134gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n644_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n848_), .A2(new_n203_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1343gat));
  INV_X1    g661(.A(new_n831_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n652_), .A2(new_n745_), .A3(new_n396_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n277_), .A3(new_n506_), .A4(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT125), .B(G141gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1344gat));
  NOR2_X1   g666(.A1(new_n831_), .A2(new_n481_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n864_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G148gat), .B1(new_n869_), .B2(new_n591_), .ZN(new_n870_));
  INV_X1    g669(.A(G148gat), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n868_), .A2(new_n871_), .A3(new_n590_), .A4(new_n864_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1345gat));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n869_), .B2(new_n635_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n868_), .A2(new_n634_), .A3(new_n864_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(new_n620_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G162gat), .B1(new_n869_), .B2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n644_), .A2(G162gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n868_), .A2(new_n864_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n652_), .A2(new_n336_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n667_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n506_), .B(new_n885_), .C1(new_n842_), .C2(new_n785_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT62), .B1(new_n886_), .B2(KEYINPUT22), .ZN(new_n887_));
  OAI21_X1  g686(.A(G169gat), .B1(new_n886_), .B2(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n234_), .B2(new_n887_), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n842_), .A2(new_n785_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n885_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G176gat), .B1(new_n893_), .B2(new_n590_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n831_), .A2(new_n667_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n591_), .A2(new_n884_), .A3(new_n235_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1349gat));
  NAND4_X1  g696(.A1(new_n895_), .A2(new_n652_), .A3(new_n336_), .A4(new_n634_), .ZN(new_n898_));
  INV_X1    g697(.A(G183gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n635_), .A2(new_n222_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n899_), .B1(new_n893_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n893_), .A2(new_n402_), .A3(new_n860_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n891_), .A2(new_n879_), .A3(new_n892_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n223_), .B2(new_n903_), .ZN(G1351gat));
  NAND2_X1  g703(.A1(new_n652_), .A2(new_n448_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n863_), .A2(new_n277_), .A3(new_n506_), .A4(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT126), .B(G197gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1352gat));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n831_), .A2(new_n481_), .A3(new_n591_), .A4(new_n905_), .ZN(new_n911_));
  INV_X1    g710(.A(G204gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n863_), .A2(new_n277_), .A3(new_n590_), .A4(new_n906_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(KEYINPUT127), .A3(G204gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n349_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n915_), .A3(new_n917_), .ZN(G1353gat));
  XNOR2_X1  g717(.A(KEYINPUT63), .B(G211gat), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n868_), .A2(new_n634_), .A3(new_n906_), .A4(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n863_), .A2(new_n277_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n921_), .A2(new_n635_), .A3(new_n905_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  NAND4_X1  g723(.A1(new_n868_), .A2(new_n340_), .A3(new_n860_), .A4(new_n906_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n921_), .A2(new_n879_), .A3(new_n905_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n340_), .ZN(G1355gat));
endmodule


