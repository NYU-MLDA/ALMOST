//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT64), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n207_), .A2(new_n209_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n208_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT7), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n221_), .C1(G99gat), .C2(G106gat), .ZN(new_n222_));
  OAI22_X1  g021(.A1(new_n220_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  AOI211_X1 g025(.A(KEYINPUT8), .B(new_n217_), .C1(new_n226_), .C2(new_n214_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n223_), .B(new_n221_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n213_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT6), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT6), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(KEYINPUT6), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n213_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n208_), .B1(new_n228_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT67), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n241_), .B(new_n208_), .C1(new_n228_), .C2(new_n238_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(KEYINPUT8), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n227_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n240_), .A2(new_n242_), .A3(KEYINPUT68), .A4(KEYINPUT8), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n216_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G57gat), .B(G64gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT69), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G78gat), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(KEYINPUT11), .A3(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n235_), .A2(new_n236_), .A3(new_n213_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n213_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n217_), .B1(new_n259_), .B2(new_n226_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT8), .B1(new_n260_), .B2(new_n241_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n242_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n244_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n227_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n246_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n215_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n255_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n256_), .A2(new_n268_), .A3(KEYINPUT12), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n255_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n203_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n202_), .B1(new_n256_), .B2(new_n268_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G176gat), .B(G204gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n273_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT13), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT34), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT35), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT15), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G29gat), .B(G36gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G43gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(G50gat), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(G50gat), .B1(new_n290_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n285_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n288_), .B(new_n289_), .ZN(new_n296_));
  INV_X1    g095(.A(G50gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(KEYINPUT15), .A3(new_n292_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n284_), .B1(new_n266_), .B2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n293_), .A2(new_n294_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT72), .B1(new_n247_), .B2(new_n302_), .ZN(new_n303_));
  AND4_X1   g102(.A1(KEYINPUT72), .A2(new_n265_), .A3(new_n215_), .A4(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n301_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n283_), .A2(KEYINPUT35), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n301_), .B(new_n306_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT73), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT36), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .A4(new_n317_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n316_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT36), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT37), .B1(new_n321_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n329_), .B(new_n326_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G231gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n255_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G1gat), .ZN(new_n334_));
  INV_X1    g133(.A(G8gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT14), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G15gat), .B(G22gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n337_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT76), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G8gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n333_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT17), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G155gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT16), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n347_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(KEYINPUT17), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n331_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n281_), .A2(new_n358_), .A3(KEYINPUT77), .ZN(new_n359_));
  AND3_X1   g158(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT22), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G169gat), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n363_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n362_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n364_), .A2(new_n368_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(KEYINPUT24), .A3(new_n371_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT26), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(KEYINPUT26), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(KEYINPUT81), .B2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n377_), .B(new_n379_), .C1(new_n385_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n374_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT30), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT31), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n393_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT84), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n402_), .B(KEYINPUT83), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n401_), .B(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G127gat), .B(G134gat), .Z(new_n405_));
  XOR2_X1   g204(.A(G113gat), .B(G120gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n404_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n398_), .A2(new_n399_), .A3(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  INV_X1    g215(.A(G155gat), .ZN(new_n417_));
  INV_X1    g216(.A(G162gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT1), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n419_), .A2(new_n421_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G141gat), .B(G148gat), .Z(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n424_), .A3(new_n420_), .ZN(new_n428_));
  INV_X1    g227(.A(G141gat), .ZN(new_n429_));
  INV_X1    g228(.A(G148gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT3), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n428_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n415_), .B1(new_n427_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n426_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT86), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G22gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n297_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT28), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G22gat), .A2(G50gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT87), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n450_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n445_), .A2(new_n458_), .ZN(new_n459_));
  AOI211_X1 g258(.A(KEYINPUT29), .B(new_n457_), .C1(new_n439_), .C2(new_n444_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n414_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n445_), .A2(new_n458_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n463_), .A2(new_n460_), .A3(KEYINPUT88), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n439_), .A2(KEYINPUT29), .A3(new_n444_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G228gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G211gat), .B(G218gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT89), .ZN(new_n469_));
  OR2_X1    g268(.A1(G197gat), .A2(G204gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G197gat), .A2(G204gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT21), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT21), .B1(new_n470_), .B2(new_n471_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G211gat), .B(G218gat), .Z(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n469_), .B(new_n472_), .C1(new_n475_), .C2(new_n474_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(new_n467_), .A3(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n440_), .A2(new_n441_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n478_), .ZN(new_n484_));
  OAI211_X1 g283(.A(G228gat), .B(G233gat), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G78gat), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n480_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n205_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n480_), .A2(new_n485_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G78gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(G106gat), .A3(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n465_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n493_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n465_), .A2(new_n489_), .A3(new_n493_), .A4(KEYINPUT90), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G29gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G85gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n439_), .A2(new_n408_), .A3(new_n444_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT94), .B1(new_n407_), .B2(new_n481_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n439_), .A2(new_n408_), .A3(KEYINPUT94), .A4(new_n444_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT4), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n439_), .A2(new_n408_), .A3(new_n513_), .A4(new_n444_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n511_), .A2(new_n512_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n513_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT95), .B1(new_n520_), .B2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n515_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n505_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n505_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT99), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n519_), .A2(new_n521_), .B1(new_n510_), .B2(new_n515_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n529_), .B(new_n530_), .C1(new_n505_), .C2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G8gat), .B(G36gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT18), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G92gat), .ZN(new_n536_));
  INV_X1    g335(.A(G64gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n534_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n211_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n390_), .A2(new_n479_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G226gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT19), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n381_), .A2(G190gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT91), .B1(new_n387_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n382_), .A2(new_n384_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n386_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n362_), .B2(new_n376_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G183gat), .A2(G190gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n555_));
  AND4_X1   g354(.A1(new_n550_), .A2(new_n376_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n549_), .B(new_n379_), .C1(new_n551_), .C2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n363_), .A2(new_n371_), .A3(new_n369_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n484_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n541_), .A2(KEYINPUT20), .A3(new_n544_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n558_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n479_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n484_), .A2(new_n374_), .A3(new_n389_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n544_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n560_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AOI211_X1 g366(.A(KEYINPUT93), .B(new_n544_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n540_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n479_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT20), .A3(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n543_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT93), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n565_), .A2(new_n566_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n540_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n560_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT27), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n541_), .A2(KEYINPUT20), .A3(new_n559_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n543_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n563_), .A2(new_n544_), .A3(new_n564_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n582_), .B2(new_n540_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n577_), .A2(new_n578_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n584_));
  AND4_X1   g383(.A1(new_n500_), .A2(new_n527_), .A3(new_n532_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT33), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n505_), .B1(new_n510_), .B2(new_n516_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n514_), .A2(new_n515_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n520_), .B2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n569_), .A2(new_n576_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n526_), .A2(new_n588_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n536_), .A2(new_n539_), .A3(KEYINPUT32), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n582_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n582_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n573_), .A2(new_n574_), .A3(new_n560_), .A4(new_n598_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n603_), .B(new_n604_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n500_), .B1(new_n596_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n413_), .B1(new_n585_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT100), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n411_), .A2(new_n412_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n587_), .B(new_n525_), .C1(new_n521_), .C2(new_n519_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n569_), .A2(new_n576_), .A3(new_n593_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(new_n589_), .A3(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT98), .B(new_n598_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n604_), .B1(new_n600_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n512_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n520_), .A2(KEYINPUT95), .A3(new_n517_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n523_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n505_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n615_), .B1(new_n620_), .B2(new_n529_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n610_), .B1(new_n613_), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n500_), .A2(new_n527_), .A3(new_n532_), .A4(new_n584_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n609_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n413_), .A2(new_n500_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n527_), .A2(new_n532_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n584_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n608_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n300_), .A2(new_n344_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT79), .Z(new_n632_));
  INV_X1    g431(.A(new_n302_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n344_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n344_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT78), .B1(new_n640_), .B2(new_n634_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n634_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT78), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n636_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n638_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT80), .ZN(new_n649_));
  XOR2_X1   g448(.A(G113gat), .B(G141gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n647_), .B(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n359_), .A2(new_n630_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT77), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n281_), .A2(new_n358_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT101), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT101), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n628_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n662_));
  INV_X1    g461(.A(new_n652_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n280_), .A2(new_n357_), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n629_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT100), .B(new_n609_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n321_), .A2(new_n327_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n628_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n661_), .A2(new_n662_), .A3(new_n671_), .ZN(G1324gat));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  INV_X1    g472(.A(new_n584_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n657_), .A2(new_n335_), .A3(new_n674_), .A4(new_n658_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n664_), .A2(new_n669_), .A3(new_n674_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n335_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT103), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT104), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n678_), .A2(new_n684_), .A3(new_n679_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n682_), .A2(KEYINPUT104), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n681_), .A2(new_n683_), .A3(new_n685_), .A4(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n675_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n683_), .B1(new_n681_), .B2(new_n685_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n673_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(KEYINPUT40), .A3(new_n675_), .A4(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n670_), .B2(new_n413_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT41), .Z(new_n695_));
  OR2_X1    g494(.A1(new_n413_), .A2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n659_), .B2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n670_), .B2(new_n610_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n500_), .A2(new_n446_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n659_), .B2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n357_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n280_), .A2(new_n702_), .A3(new_n663_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n668_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n667_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n628_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(new_n328_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n330_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n630_), .B2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n608_), .A2(new_n626_), .A3(KEYINPUT105), .A4(new_n629_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n711_), .A2(new_n712_), .A3(new_n710_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n667_), .B2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n328_), .A2(new_n330_), .A3(KEYINPUT43), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n630_), .A2(new_n721_), .A3(KEYINPUT106), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n703_), .C1(new_n717_), .C2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(G29gat), .A3(new_n708_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n630_), .A2(new_n721_), .A3(KEYINPUT106), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT106), .B1(new_n630_), .B2(new_n721_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n714_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n331_), .A3(new_n716_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT43), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT44), .B1(new_n732_), .B2(new_n703_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n709_), .B1(new_n725_), .B2(new_n734_), .ZN(G1328gat));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n584_), .A2(G36gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OR3_X1    g538(.A1(new_n706_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n706_), .B2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n724_), .A2(new_n674_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G36gat), .B1(new_n743_), .B2(new_n733_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(KEYINPUT107), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(G36gat), .C1(new_n743_), .C2(new_n733_), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT109), .B(new_n736_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(KEYINPUT107), .ZN(new_n749_));
  INV_X1    g548(.A(new_n742_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n747_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n748_), .A2(new_n753_), .ZN(G1329gat));
  OAI21_X1  g553(.A(new_n289_), .B1(new_n706_), .B2(new_n413_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n724_), .A2(G43gat), .A3(new_n609_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n733_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT110), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT110), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(KEYINPUT47), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT47), .B1(new_n758_), .B2(new_n759_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1330gat));
  NAND3_X1  g561(.A1(new_n707_), .A2(new_n297_), .A3(new_n500_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n724_), .A2(new_n500_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n733_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G50gat), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n765_), .A2(new_n733_), .A3(new_n764_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT112), .ZN(G1331gat));
  NOR2_X1   g569(.A1(new_n281_), .A2(new_n652_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n702_), .A3(new_n669_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G57gat), .B1(new_n772_), .B2(new_n628_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n358_), .A3(new_n630_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n628_), .A2(G57gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(G1332gat));
  OAI21_X1  g575(.A(G64gat), .B1(new_n772_), .B2(new_n584_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT48), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n674_), .A2(new_n537_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n774_), .B2(new_n779_), .ZN(G1333gat));
  OR3_X1    g579(.A1(new_n774_), .A2(G71gat), .A3(new_n413_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G71gat), .B1(new_n772_), .B2(new_n413_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(KEYINPUT113), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(KEYINPUT113), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(KEYINPUT49), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT49), .B1(new_n784_), .B2(new_n785_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  OAI21_X1  g587(.A(G78gat), .B1(new_n772_), .B2(new_n610_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT50), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n500_), .A2(new_n486_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT114), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n774_), .B2(new_n792_), .ZN(G1335gat));
  NOR3_X1   g592(.A1(new_n281_), .A2(new_n702_), .A3(new_n652_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n705_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT115), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n210_), .A3(new_n708_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n732_), .A2(new_n794_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n708_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(new_n210_), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n211_), .A3(new_n674_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n798_), .A2(new_n674_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n211_), .ZN(G1337gat));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n609_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n609_), .A2(new_n204_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n804_), .A2(G99gat), .B1(new_n796_), .B2(new_n805_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g606(.A1(new_n796_), .A2(new_n205_), .A3(new_n500_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n798_), .A2(new_n500_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(G106gat), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT52), .B(new_n205_), .C1(new_n798_), .C2(new_n500_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT53), .ZN(G1339gat));
  OR3_X1    g613(.A1(new_n655_), .A2(KEYINPUT54), .A3(new_n652_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n655_), .B2(new_n652_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n632_), .A2(new_n642_), .A3(new_n636_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n651_), .B1(new_n645_), .B2(new_n635_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n638_), .A2(new_n646_), .A3(new_n651_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n278_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n273_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n819_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n273_), .A2(new_n825_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT119), .A3(new_n823_), .A4(new_n822_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n269_), .A2(new_n270_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT55), .B1(new_n831_), .B2(new_n202_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n271_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n271_), .A2(new_n835_), .A3(KEYINPUT55), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n202_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT116), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n825_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n833_), .A2(new_n832_), .B1(new_n837_), .B2(KEYINPUT116), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n278_), .B1(new_n843_), .B2(new_n836_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(KEYINPUT56), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n830_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n830_), .B(KEYINPUT58), .C1(new_n842_), .C2(new_n845_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(new_n331_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n841_), .B1(new_n844_), .B2(KEYINPUT117), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n840_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n851_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n853_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n844_), .A2(KEYINPUT117), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(KEYINPUT118), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n842_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n855_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n663_), .A2(new_n826_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n279_), .A2(new_n824_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n668_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n850_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n863_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n668_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n818_), .B1(new_n871_), .B2(new_n357_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n627_), .A2(new_n708_), .A3(new_n584_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n865_), .B2(new_n704_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n848_), .A2(new_n331_), .A3(new_n849_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n867_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n869_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n357_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n817_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  INV_X1    g680(.A(new_n873_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n883_), .A3(new_n652_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G113gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n872_), .A2(new_n873_), .ZN(new_n886_));
  INV_X1    g685(.A(G113gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n652_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1340gat));
  NAND3_X1  g688(.A1(new_n874_), .A2(new_n883_), .A3(new_n280_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(G120gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n886_), .B(new_n894_), .C1(KEYINPUT60), .C2(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1341gat));
  NAND3_X1  g695(.A1(new_n874_), .A2(new_n883_), .A3(new_n702_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G127gat), .ZN(new_n898_));
  INV_X1    g697(.A(G127gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n886_), .A2(new_n899_), .A3(new_n702_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1342gat));
  AND2_X1   g700(.A1(new_n874_), .A2(new_n883_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT122), .B(G134gat), .Z(new_n903_));
  NOR2_X1   g702(.A1(new_n713_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n702_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n668_), .B(new_n882_), .C1(new_n905_), .C2(new_n818_), .ZN(new_n906_));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT121), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n910_), .A3(new_n907_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n902_), .A2(new_n904_), .B1(new_n909_), .B2(new_n911_), .ZN(G1343gat));
  NOR2_X1   g711(.A1(new_n610_), .A2(new_n609_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n628_), .A2(new_n674_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n913_), .B(new_n914_), .C1(new_n905_), .C2(new_n818_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n663_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n429_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n281_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n430_), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n915_), .A2(new_n357_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT61), .B(G155gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n915_), .B2(new_n713_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n668_), .A2(new_n418_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n915_), .B2(new_n924_), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n708_), .A2(new_n413_), .A3(new_n584_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n652_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT123), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n880_), .A2(new_n610_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(new_n930_), .A3(G169gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n880_), .A2(new_n610_), .A3(new_n926_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n652_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n931_), .A2(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1348gat));
  OAI21_X1  g734(.A(new_n368_), .B1(new_n933_), .B2(new_n281_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n872_), .A2(new_n500_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n937_), .A2(G176gat), .A3(new_n280_), .A4(new_n926_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n933_), .A2(new_n357_), .A3(new_n386_), .ZN(new_n940_));
  INV_X1    g739(.A(G183gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n937_), .A2(new_n702_), .A3(new_n926_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n933_), .B2(new_n713_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n668_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n933_), .B2(new_n945_), .ZN(G1351gat));
  NAND3_X1  g745(.A1(new_n913_), .A2(new_n628_), .A3(new_n674_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n879_), .B2(new_n817_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n652_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n280_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT124), .B(G204gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1353gat));
  INV_X1    g752(.A(new_n947_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n357_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n955_), .B(KEYINPUT125), .Z(new_n956_));
  OAI211_X1 g755(.A(new_n954_), .B(new_n956_), .C1(new_n905_), .C2(new_n818_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(KEYINPUT126), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n880_), .A2(new_n960_), .A3(new_n954_), .A4(new_n956_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n958_), .A2(new_n959_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n958_), .B2(new_n961_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1354gat));
  AOI21_X1  g763(.A(new_n315_), .B1(new_n948_), .B2(new_n331_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n704_), .A2(G218gat), .ZN(new_n966_));
  AND3_X1   g765(.A1(new_n880_), .A2(new_n954_), .A3(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(new_n965_), .B2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n948_), .A2(new_n966_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n872_), .A2(new_n713_), .A3(new_n947_), .ZN(new_n971_));
  OAI211_X1 g770(.A(new_n969_), .B(new_n970_), .C1(new_n971_), .C2(new_n315_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n968_), .A2(new_n972_), .ZN(G1355gat));
endmodule


