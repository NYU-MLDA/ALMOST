//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n208_), .B(new_n209_), .Z(new_n210_));
  XNOR2_X1  g009(.A(G71gat), .B(G78gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n211_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n210_), .B(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G155gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G183gat), .B(G211gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT17), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n218_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n225_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(KEYINPUT76), .Z(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G190gat), .B(G218gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G134gat), .B(G162gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT36), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT35), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n241_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT73), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT6), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT66), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G85gat), .B(G92gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT8), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n253_), .A2(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT10), .B(G99gat), .Z(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  AOI22_X1  g064(.A1(KEYINPUT9), .A2(new_n256_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n266_), .B(new_n251_), .C1(KEYINPUT9), .C2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT65), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G43gat), .B(G50gat), .ZN(new_n271_));
  INV_X1    g070(.A(G36gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT70), .B(G29gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n275_), .B(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n245_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n268_), .B(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n261_), .B1(new_n257_), .B2(KEYINPUT8), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n263_), .A2(new_n269_), .A3(KEYINPUT67), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n275_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n281_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n279_), .A2(new_n280_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n243_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n243_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n294_), .A2(new_n279_), .A3(new_n245_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n237_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n236_), .A2(KEYINPUT36), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT37), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT37), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(KEYINPUT24), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT25), .B(G183gat), .Z(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n312_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT82), .B1(new_n312_), .B2(KEYINPUT23), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n315_), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n305_), .A2(KEYINPUT24), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT94), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n314_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(G183gat), .A3(G190gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT94), .ZN(new_n324_));
  INV_X1    g123(.A(new_n318_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n311_), .B1(new_n319_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n312_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT80), .B1(new_n312_), .B2(KEYINPUT23), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n321_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n315_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n328_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  AOI211_X1 g138(.A(KEYINPUT96), .B(new_n337_), .C1(new_n331_), .C2(new_n335_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT95), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n306_), .B1(new_n343_), .B2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n327_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  INV_X1    g146(.A(G218gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT90), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT90), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(G218gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(G211gat), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(G218gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(KEYINPUT90), .ZN(new_n354_));
  INV_X1    g153(.A(G211gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n347_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  INV_X1    g157(.A(G204gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G197gat), .ZN(new_n360_));
  INV_X1    g159(.A(G197gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G204gat), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n357_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n358_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n355_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT89), .B(new_n365_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n363_), .A2(new_n358_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT97), .B1(new_n346_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n369_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n357_), .A3(new_n365_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n369_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT91), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G183gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT78), .B(G183gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT79), .B1(new_n382_), .B2(KEYINPUT25), .ZN(new_n385_));
  OAI221_X1 g184(.A(new_n308_), .B1(KEYINPUT25), .B2(new_n381_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n336_), .A2(new_n325_), .A3(new_n307_), .ZN(new_n387_));
  INV_X1    g186(.A(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n323_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n306_), .ZN(new_n391_));
  INV_X1    g190(.A(G176gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n342_), .B2(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n386_), .A2(new_n387_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n373_), .B1(new_n380_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n371_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT97), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n344_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n397_), .C1(new_n398_), .C2(new_n327_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n372_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n373_), .B1(new_n346_), .B2(new_n371_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n394_), .B2(new_n380_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(new_n403_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n400_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n412_));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n406_), .A2(new_n409_), .A3(new_n418_), .A4(new_n410_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT106), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n408_), .A2(new_n403_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n403_), .B2(new_n400_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n416_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n425_), .B2(KEYINPUT105), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n419_), .C1(KEYINPUT105), .C2(new_n425_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT1), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G155gat), .A3(G162gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT86), .ZN(new_n441_));
  NOR3_X1   g240(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT3), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n436_), .B(KEYINPUT2), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT28), .B1(new_n447_), .B2(KEYINPUT29), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n440_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n431_), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n429_), .B(new_n451_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT28), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G22gat), .B(G50gat), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n448_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n396_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(G228gat), .A3(G233gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n380_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n447_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT88), .B1(new_n447_), .B2(KEYINPUT29), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n463_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT92), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n469_), .B2(new_n460_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n472_));
  OR3_X1    g271(.A1(new_n460_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G78gat), .B(G106gat), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n428_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G127gat), .B(G134gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G120gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n441_), .A2(new_n486_), .A3(new_n446_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT101), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT101), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n453_), .A2(new_n491_), .A3(new_n486_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n483_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n488_), .A2(KEYINPUT4), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(KEYINPUT4), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n496_), .B2(new_n483_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(G85gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT103), .B1(new_n498_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(KEYINPUT103), .A3(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n486_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G15gat), .B(G43gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT84), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n511_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(new_n394_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G71gat), .B(G99gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n515_), .B(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n509_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n481_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n400_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT98), .B1(new_n400_), .B2(new_n403_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n418_), .B1(new_n527_), .B2(new_n409_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n419_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT100), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n496_), .A2(new_n482_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n503_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n482_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT33), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n496_), .A2(new_n483_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n493_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(KEYINPUT33), .A3(new_n536_), .A4(new_n502_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT102), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n497_), .A2(KEYINPUT102), .A3(KEYINPUT33), .A4(new_n502_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n534_), .A2(new_n505_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT100), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n417_), .A2(new_n542_), .A3(new_n419_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n530_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n411_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n424_), .A2(new_n545_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n506_), .A2(new_n546_), .A3(new_n507_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n480_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT104), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT104), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n552_), .A3(new_n480_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n421_), .A2(new_n508_), .A3(new_n479_), .A4(new_n427_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n521_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n524_), .B1(new_n556_), .B2(KEYINPUT107), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT107), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n558_), .A3(new_n521_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n232_), .B(new_n304_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT64), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n288_), .A2(new_n217_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n288_), .A2(new_n217_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n217_), .B(new_n226_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n288_), .A2(new_n217_), .B1(new_n568_), .B2(KEYINPUT12), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n288_), .B2(new_n217_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n571_), .A3(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT5), .B(G176gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n572_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n275_), .B(new_n208_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n586_), .A2(KEYINPUT77), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT77), .B1(new_n586_), .B2(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n587_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n289_), .A2(new_n277_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n586_), .B2(new_n277_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n588_), .B(new_n589_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n593_), .B(new_n596_), .Z(new_n597_));
  NOR2_X1   g396(.A1(new_n585_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n560_), .A2(new_n203_), .A3(new_n509_), .A4(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT108), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n420_), .A2(KEYINPUT106), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT106), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n604_), .B(KEYINPUT27), .C1(new_n417_), .C2(new_n419_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n479_), .B(new_n427_), .C1(new_n603_), .C2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n509_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n552_), .B1(new_n549_), .B2(new_n480_), .ZN(new_n608_));
  AOI211_X1 g407(.A(KEYINPUT104), .B(new_n479_), .C1(new_n544_), .C2(new_n548_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n521_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT107), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n524_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n559_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n300_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n598_), .A2(new_n231_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT109), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n509_), .A3(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n601_), .A2(new_n599_), .B1(new_n620_), .B2(G1gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n600_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n602_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT110), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1324gat));
  AND2_X1   g424(.A1(new_n560_), .A2(new_n598_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n428_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n204_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n627_), .A3(new_n619_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n629_), .B2(G8gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n617_), .A2(new_n619_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n611_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n626_), .A2(new_n636_), .A3(new_n611_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n637_), .B2(new_n479_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n626_), .A2(new_n642_), .A3(new_n479_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n598_), .A2(new_n232_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n615_), .A2(new_n300_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n509_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n647_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT111), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n304_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n652_), .B1(new_n614_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n304_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n651_), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(new_n651_), .C1(new_n656_), .C2(new_n660_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n508_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n650_), .B1(new_n666_), .B2(new_n649_), .ZN(G1328gat));
  NOR2_X1   g466(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n668_));
  INV_X1    g467(.A(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n614_), .A2(new_n658_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n654_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n652_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(new_n651_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n627_), .B1(new_n669_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n614_), .A2(new_n616_), .A3(new_n651_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(G36gat), .A3(new_n428_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n668_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n428_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n668_), .B(new_n680_), .C1(new_n682_), .C2(new_n272_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1329gat));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n611_), .B1(new_n669_), .B2(new_n674_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G43gat), .ZN(new_n688_));
  INV_X1    g487(.A(G43gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n648_), .A2(new_n689_), .A3(new_n611_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n686_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n521_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n686_), .B(new_n690_), .C1(new_n692_), .C2(new_n689_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n648_), .A2(new_n696_), .A3(new_n479_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n480_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n696_), .ZN(G1331gat));
  INV_X1    g498(.A(new_n585_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n597_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n617_), .A2(new_n231_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n508_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n560_), .A2(new_n702_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n509_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n703_), .B2(new_n428_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  INV_X1    g509(.A(G64gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n711_), .A3(new_n627_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1333gat));
  OAI21_X1  g512(.A(G71gat), .B1(new_n703_), .B2(new_n521_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n716_), .A3(new_n611_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n703_), .B2(new_n480_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n721_), .A3(new_n479_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n702_), .A2(new_n232_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n615_), .A2(new_n300_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(G85gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n509_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n724_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n673_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n508_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n727_), .B1(new_n733_), .B2(new_n726_), .ZN(G1336gat));
  INV_X1    g533(.A(G92gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n735_), .A3(new_n627_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n428_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n735_), .ZN(G1337gat));
  NAND3_X1  g537(.A1(new_n673_), .A2(new_n611_), .A3(new_n728_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G99gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n725_), .A2(new_n264_), .A3(new_n611_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g542(.A1(new_n725_), .A2(new_n265_), .A3(new_n479_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n479_), .B(new_n728_), .C1(new_n656_), .C2(new_n660_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT54), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT54), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n302_), .A2(new_n597_), .A3(new_n231_), .A4(new_n303_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n752_), .B(new_n753_), .C1(new_n754_), .C2(new_n585_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n585_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n753_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n562_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n572_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT55), .A4(new_n562_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n577_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n579_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT117), .B1(new_n769_), .B2(new_n766_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n701_), .A2(new_n580_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n593_), .A2(new_n596_), .ZN(new_n774_));
  MUX2_X1   g573(.A(new_n586_), .B(new_n592_), .S(new_n590_), .Z(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n596_), .B2(new_n775_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n772_), .A2(new_n773_), .B1(new_n581_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n758_), .B1(new_n777_), .B2(new_n616_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n777_), .A2(new_n758_), .A3(new_n616_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n776_), .A2(new_n580_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n786_));
  INV_X1    g585(.A(new_n770_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n785_), .B(KEYINPUT58), .C1(new_n787_), .C2(new_n786_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n304_), .A3(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT118), .B(new_n758_), .C1(new_n777_), .C2(new_n616_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n780_), .A2(new_n782_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n757_), .B1(new_n794_), .B2(new_n232_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n481_), .A2(new_n508_), .A3(new_n521_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n795_), .A2(KEYINPUT120), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT120), .B1(new_n795_), .B2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n701_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n792_), .A2(new_n778_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n781_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n792_), .A2(new_n778_), .A3(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n757_), .B1(new_n806_), .B2(new_n232_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n797_), .A2(KEYINPUT59), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT122), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n797_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n231_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n812_), .B(new_n808_), .C1(new_n813_), .C2(new_n757_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n810_), .A2(KEYINPUT123), .A3(new_n811_), .A4(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n597_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n801_), .B1(new_n819_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n815_), .B2(new_n700_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT60), .ZN(new_n822_));
  AOI21_X1  g621(.A(G120gat), .B1(new_n585_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(G120gat), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(KEYINPUT124), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT124), .B1(new_n824_), .B2(new_n825_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n826_), .B2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n800_), .B2(new_n231_), .ZN(new_n829_));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(new_n231_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n800_), .B2(new_n616_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n657_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g634(.A1(new_n795_), .A2(new_n611_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n606_), .A2(new_n508_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n597_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n437_), .ZN(G1344gat));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n700_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n438_), .ZN(G1345gat));
  OR3_X1    g641(.A1(new_n838_), .A2(KEYINPUT125), .A3(new_n232_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT125), .B1(new_n838_), .B2(new_n232_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(new_n838_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n849_), .A2(G162gat), .A3(new_n655_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G162gat), .B1(new_n849_), .B2(new_n616_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  INV_X1    g651(.A(new_n807_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n428_), .A2(new_n479_), .A3(new_n523_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G169gat), .B1(new_n855_), .B2(new_n597_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n856_), .A2(KEYINPUT62), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(KEYINPUT62), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n597_), .A2(new_n343_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT126), .Z(new_n860_));
  OAI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n855_), .B2(new_n860_), .ZN(G1348gat));
  INV_X1    g660(.A(new_n855_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G176gat), .B1(new_n862_), .B2(new_n585_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n795_), .A2(new_n479_), .A3(new_n428_), .A4(new_n523_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n700_), .A2(new_n392_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  AND2_X1   g665(.A1(new_n231_), .A2(new_n310_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n231_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n862_), .A2(new_n867_), .B1(new_n868_), .B2(new_n382_), .ZN(G1350gat));
  NAND3_X1  g668(.A1(new_n862_), .A2(new_n616_), .A3(new_n308_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G190gat), .B1(new_n855_), .B2(new_n657_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1351gat));
  NOR2_X1   g671(.A1(new_n480_), .A2(new_n509_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n795_), .A2(new_n611_), .A3(new_n428_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n701_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n585_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n875_), .A2(new_n231_), .A3(new_n880_), .A4(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(KEYINPUT127), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(KEYINPUT127), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n875_), .B2(new_n231_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(G1354gat));
  AOI21_X1  g685(.A(G218gat), .B1(new_n875_), .B2(new_n616_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n875_), .A2(new_n304_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(G218gat), .B2(new_n888_), .ZN(G1355gat));
endmodule


