//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  OR2_X1    g000(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n202_));
  AND2_X1   g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n202_), .A2(new_n203_), .A3(new_n206_), .A4(new_n204_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT85), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT22), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G169gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT25), .B1(new_n210_), .B2(KEYINPUT82), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G190gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n219_), .A2(new_n215_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OR3_X1    g036(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n203_), .B1(new_n202_), .B2(new_n204_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n240_));
  OAI211_X1 g039(.A(KEYINPUT84), .B(new_n238_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n204_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n207_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n240_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT84), .B1(new_n247_), .B2(new_n238_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n226_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n249_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT87), .B(G43gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT89), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n257_), .A2(new_n262_), .A3(KEYINPUT89), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n264_), .A2(KEYINPUT31), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT31), .B1(new_n264_), .B2(new_n265_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT88), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n256_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n256_), .A2(new_n270_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G85gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G57gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT99), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n264_), .A2(new_n265_), .ZN(new_n284_));
  INV_X1    g083(.A(G141gat), .ZN(new_n285_));
  INV_X1    g084(.A(G148gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(KEYINPUT90), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT3), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT90), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n288_), .A2(new_n291_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n289_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n302_), .A2(new_n292_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n305_), .A3(new_n298_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n284_), .A2(new_n308_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n296_), .A2(new_n300_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n260_), .A2(new_n263_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n283_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT4), .B1(new_n284_), .B2(new_n308_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n280_), .B(new_n282_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n312_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n316_), .B2(KEYINPUT4), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(new_n281_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT99), .B1(new_n316_), .B2(new_n282_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n279_), .B(new_n315_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n309_), .A2(new_n312_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n280_), .B1(new_n322_), .B2(new_n281_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n281_), .B2(new_n317_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n279_), .B1(new_n324_), .B2(new_n315_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n274_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT103), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT18), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT100), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT96), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n224_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT97), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n338_), .A2(new_n223_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n338_), .B2(new_n223_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n245_), .A2(new_n246_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  AND2_X1   g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G197gat), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G218gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G211gat), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(KEYINPUT21), .A3(new_n350_), .A4(new_n351_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n209_), .A2(new_n213_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n229_), .A2(G183gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n231_), .A2(new_n233_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n238_), .A3(new_n236_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n354_), .B(new_n360_), .C1(new_n361_), .C2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n336_), .B(KEYINPUT20), .C1(new_n343_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n354_), .A2(new_n360_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n249_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n209_), .A2(new_n213_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n365_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND4_X1   g172(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n224_), .B(KEYINPUT96), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT97), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n212_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n338_), .A2(new_n223_), .A3(new_n339_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n336_), .B1(new_n380_), .B2(KEYINPUT20), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n335_), .B1(new_n370_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n240_), .B1(new_n384_), .B2(new_n207_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n235_), .A2(KEYINPUT24), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n241_), .A3(new_n237_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n368_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n226_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT20), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n371_), .A2(new_n372_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n341_), .A2(new_n342_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT98), .B1(new_n393_), .B2(new_n378_), .ZN(new_n394_));
  AND4_X1   g193(.A1(KEYINPUT98), .A2(new_n376_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n391_), .B1(new_n396_), .B2(new_n368_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n335_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n382_), .A2(KEYINPUT101), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT101), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n335_), .C1(new_n370_), .C2(new_n381_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n333_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n335_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n369_), .B(new_n404_), .C1(new_n396_), .C2(new_n368_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(new_n333_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT27), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n329_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n333_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n396_), .A2(new_n368_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n391_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n398_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n389_), .B1(new_n388_), .B2(new_n226_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n403_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n336_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n366_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT100), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n398_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n412_), .B1(new_n418_), .B2(new_n400_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n401_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n406_), .A2(KEYINPUT27), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT103), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n408_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n310_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(G228gat), .A2(G233gat), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n426_), .A2(new_n389_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n310_), .B2(new_n425_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n294_), .A2(new_n295_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n290_), .B1(new_n289_), .B2(KEYINPUT90), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n299_), .B1(new_n434_), .B2(new_n291_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n304_), .A2(new_n306_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT92), .B(KEYINPUT29), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n437_), .A3(new_n368_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n438_), .A2(KEYINPUT93), .A3(new_n427_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT93), .B1(new_n438_), .B2(new_n427_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n310_), .A2(new_n425_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n444_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G22gat), .B(G50gat), .Z(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n448_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n442_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n429_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n443_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n438_), .A2(new_n427_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n438_), .A2(KEYINPUT93), .A3(new_n427_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n428_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n455_), .B1(new_n460_), .B2(new_n452_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n441_), .A2(KEYINPUT95), .A3(new_n442_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n453_), .A2(KEYINPUT94), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n452_), .A4(new_n429_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n451_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n454_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n405_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n409_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT27), .B1(new_n471_), .B2(new_n406_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n424_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(KEYINPUT104), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT104), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n408_), .B2(new_n423_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(new_n469_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n328_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n467_), .A2(new_n468_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n454_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n482_), .A3(new_n326_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n484_));
  OAI22_X1  g283(.A1(new_n321_), .A2(new_n325_), .B1(new_n470_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT102), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT102), .B(new_n484_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n324_), .A2(new_n315_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT33), .A3(new_n278_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n278_), .B1(new_n322_), .B2(new_n282_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n282_), .B2(new_n317_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n325_), .A2(KEYINPUT33), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n471_), .A2(new_n406_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n469_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n483_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n274_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n479_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT79), .ZN(new_n504_));
  INV_X1    g303(.A(G22gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n251_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G15gat), .A2(G22gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G1gat), .A2(G8gat), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n506_), .A2(new_n507_), .B1(KEYINPUT14), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n504_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G29gat), .B(G36gat), .Z(new_n511_));
  XOR2_X1   g310(.A(G43gat), .B(G50gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n510_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n513_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n510_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n515_), .A2(new_n517_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G113gat), .B(G141gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n522_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n502_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT6), .ZN(new_n532_));
  OAI22_X1  g331(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n533_));
  OR4_X1    g332(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G85gat), .ZN(new_n536_));
  INV_X1    g335(.A(G92gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT68), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT68), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n529_), .B(new_n530_), .C1(new_n535_), .C2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n532_), .A2(new_n534_), .A3(new_n533_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n528_), .A3(KEYINPUT8), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT9), .ZN(new_n549_));
  INV_X1    g348(.A(new_n539_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n538_), .C1(new_n550_), .C2(KEYINPUT66), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n532_), .A2(new_n551_), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n540_), .A2(KEYINPUT66), .A3(new_n549_), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT10), .B(G99gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT64), .B(G106gat), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n554_), .A2(KEYINPUT65), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT65), .B1(new_n554_), .B2(new_n555_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n552_), .B(new_n553_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n545_), .A2(new_n548_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n561_), .A2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n559_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT70), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n545_), .A2(new_n548_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n558_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n568_), .A2(KEYINPUT12), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT12), .B1(new_n559_), .B2(new_n568_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n559_), .A2(new_n568_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n583_), .A3(new_n570_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n569_), .A2(new_n585_), .A3(new_n571_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT73), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n573_), .A2(new_n584_), .A3(new_n586_), .A4(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n587_), .A2(KEYINPUT74), .A3(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT75), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(KEYINPUT75), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n598_), .A2(KEYINPUT75), .A3(new_n601_), .A4(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT34), .Z(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT76), .B(KEYINPUT35), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n559_), .B2(new_n514_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n577_), .B2(new_n520_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT77), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT36), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n623_), .B(KEYINPUT36), .Z(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT78), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n608_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n625_), .A2(KEYINPUT78), .A3(KEYINPUT37), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n567_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(new_n510_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT81), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(G183gat), .B(G211gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n635_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n632_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n607_), .A2(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n527_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n326_), .A2(G1gat), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n328_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n474_), .A2(KEYINPUT104), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n477_), .A2(new_n476_), .A3(new_n469_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n273_), .B1(new_n483_), .B2(new_n499_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n628_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n526_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n606_), .A2(new_n662_), .A3(new_n647_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n326_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n651_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n653_), .A2(new_n665_), .A3(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(new_n477_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n668_), .A3(new_n663_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(G8gat), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n669_), .B2(G8gat), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n477_), .A2(G8gat), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n672_), .A2(new_n673_), .B1(new_n650_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n675_), .B(new_n676_), .Z(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n664_), .B2(new_n274_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n650_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n251_), .A3(new_n273_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n681_), .A3(new_n683_), .ZN(G1326gat));
  OAI21_X1  g483(.A(G22gat), .B1(new_n664_), .B2(new_n469_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT42), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(new_n505_), .A3(new_n482_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1327gat));
  NOR3_X1   g487(.A1(new_n606_), .A2(new_n646_), .A3(new_n628_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n502_), .A2(new_n526_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n327_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n632_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n632_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n606_), .A2(new_n662_), .A3(new_n646_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(new_n698_), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n700_), .B(new_n701_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n327_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n692_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  NOR2_X1   g504(.A1(new_n477_), .A2(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n691_), .A2(KEYINPUT45), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708_));
  INV_X1    g507(.A(new_n706_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n690_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n699_), .A2(new_n702_), .A3(new_n477_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT46), .B1(new_n715_), .B2(KEYINPUT108), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n695_), .B1(new_n502_), .B2(new_n632_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n696_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n698_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n700_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n668_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n711_), .B1(new_n722_), .B2(G36gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n716_), .A2(new_n726_), .ZN(G1329gat));
  AOI21_X1  g526(.A(G43gat), .B1(new_n691_), .B2(new_n273_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n273_), .A2(G43gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n703_), .B2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n703_), .A2(new_n482_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G50gat), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n690_), .A2(G50gat), .A3(new_n469_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT109), .B(new_n735_), .C1(new_n733_), .C2(G50gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1331gat));
  NAND2_X1  g538(.A1(new_n502_), .A2(new_n662_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n648_), .A2(new_n606_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT110), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n326_), .A2(G57gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n607_), .A2(new_n526_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n661_), .A2(new_n646_), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n326_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n477_), .A2(G64gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n747_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n751_), .B2(new_n477_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1333gat));
  NOR2_X1   g557(.A1(new_n274_), .A2(G71gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n746_), .A2(new_n747_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G71gat), .B1(new_n751_), .B2(new_n274_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n469_), .A2(G78gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n747_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G78gat), .B1(new_n751_), .B2(new_n469_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1335gat));
  AND3_X1   g567(.A1(new_n697_), .A2(new_n647_), .A3(new_n750_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n327_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n606_), .A2(new_n647_), .A3(new_n660_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n742_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n327_), .A2(new_n536_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(new_n770_), .A2(new_n536_), .B1(new_n773_), .B2(new_n774_), .ZN(G1336gat));
  AND2_X1   g574(.A1(new_n769_), .A2(new_n668_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n668_), .A2(new_n537_), .ZN(new_n777_));
  OAI22_X1  g576(.A1(new_n776_), .A2(new_n537_), .B1(new_n773_), .B2(new_n777_), .ZN(G1337gat));
  NAND4_X1  g577(.A1(new_n742_), .A2(new_n273_), .A3(new_n554_), .A4(new_n772_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n769_), .A2(new_n273_), .ZN(new_n780_));
  INV_X1    g579(.A(G99gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g582(.A1(new_n697_), .A2(new_n482_), .A3(new_n647_), .A4(new_n750_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n482_), .A2(new_n555_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n786_), .A2(new_n787_), .B1(new_n773_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g589(.A(new_n525_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n521_), .B(new_n517_), .C1(new_n510_), .C2(new_n514_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n522_), .A2(new_n525_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n597_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n570_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n584_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n580_), .A2(new_n583_), .A3(KEYINPUT55), .A4(new_n570_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n594_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n593_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT114), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n799_), .A2(new_n594_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n801_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n594_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(KEYINPUT58), .A4(new_n794_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n803_), .A2(new_n804_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n805_), .A2(new_n811_), .A3(new_n632_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n526_), .A2(new_n597_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n598_), .A2(new_n599_), .A3(new_n793_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n628_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n813_), .B(new_n819_), .C1(new_n820_), .C2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n647_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n649_), .B2(new_n526_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n607_), .A2(new_n648_), .A3(new_n824_), .A4(new_n662_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n326_), .B(new_n274_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n813_), .A2(new_n819_), .A3(KEYINPUT116), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT116), .B1(new_n813_), .B2(new_n819_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n817_), .A2(new_n820_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n826_), .B1(new_n834_), .B2(new_n646_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT115), .ZN(new_n838_));
  MUX2_X1   g637(.A(KEYINPUT115), .B(new_n838_), .S(new_n828_), .Z(new_n839_));
  OAI21_X1  g638(.A(new_n830_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n662_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n662_), .A2(G113gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n829_), .B2(new_n842_), .ZN(G1340gat));
  INV_X1    g642(.A(new_n829_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n845_));
  AOI21_X1  g644(.A(G120gat), .B1(new_n606_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n845_), .B2(G120gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G120gat), .B1(new_n840_), .B2(new_n607_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n844_), .B2(new_n646_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n840_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n647_), .A2(KEYINPUT118), .ZN(new_n855_));
  MUX2_X1   g654(.A(KEYINPUT118), .B(new_n855_), .S(G127gat), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1342gat));
  AOI21_X1  g656(.A(G134gat), .B1(new_n844_), .B2(new_n660_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n632_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT119), .B(G134gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n854_), .B2(new_n861_), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n469_), .A2(new_n326_), .A3(new_n273_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n827_), .A2(new_n477_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n662_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n285_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n607_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT120), .B(G148gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1345gat));
  NOR2_X1   g668(.A1(new_n864_), .A2(new_n647_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT61), .B(G155gat), .Z(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  NAND2_X1  g671(.A1(new_n632_), .A2(G162gat), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT122), .Z(new_n874_));
  NOR2_X1   g673(.A1(new_n864_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n864_), .B2(new_n628_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n877_), .A2(KEYINPUT121), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT121), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n654_), .A2(new_n477_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n482_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n813_), .A2(new_n819_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n833_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n813_), .A2(new_n819_), .A3(KEYINPUT116), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n646_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n826_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n526_), .B(new_n883_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n835_), .A2(new_n892_), .A3(new_n526_), .A4(new_n883_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n893_), .A3(G169gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n883_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n886_), .A2(new_n887_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n647_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n826_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(new_n220_), .A3(new_n222_), .A4(new_n526_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n891_), .A2(new_n893_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n896_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  AOI22_X1  g702(.A1(new_n647_), .A2(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT124), .B1(new_n904_), .B2(new_n482_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n827_), .A2(new_n906_), .A3(new_n469_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n907_), .A3(new_n881_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n606_), .A2(G176gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n216_), .A2(new_n218_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n900_), .B2(new_n606_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT125), .B1(new_n910_), .B2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n835_), .A2(new_n606_), .A3(new_n883_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n916_), .B(new_n917_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n918_), .ZN(G1349gat));
  OR2_X1    g718(.A1(new_n908_), .A2(new_n647_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n647_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n920_), .A2(new_n210_), .B1(new_n900_), .B2(new_n921_), .ZN(G1350gat));
  INV_X1    g721(.A(new_n900_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G190gat), .B1(new_n923_), .B2(new_n859_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n660_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(new_n925_), .ZN(G1351gat));
  NOR4_X1   g725(.A1(new_n477_), .A2(new_n469_), .A3(new_n327_), .A4(new_n273_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n827_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n662_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n348_), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n607_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(G204gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1353gat));
  INV_X1    g732(.A(new_n928_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n646_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n928_), .B2(new_n859_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n660_), .A2(new_n355_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n928_), .B2(new_n941_), .ZN(G1355gat));
endmodule


