//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(KEYINPUT7), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT66), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT8), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(KEYINPUT8), .B(new_n202_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT9), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(new_n202_), .B2(KEYINPUT9), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  AND3_X1   g018(.A1(new_n219_), .A2(KEYINPUT65), .A3(new_n206_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n219_), .B2(new_n206_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n204_), .B(new_n218_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n213_), .A2(new_n214_), .A3(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n226_), .B(KEYINPUT15), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT35), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n230_), .A3(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G190gat), .B(G218gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT69), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G134gat), .B(G162gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT36), .ZN(new_n244_));
  INV_X1    g043(.A(new_n238_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n228_), .A2(new_n245_), .A3(new_n230_), .A4(new_n236_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n239_), .A2(KEYINPUT70), .A3(new_n244_), .A4(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n239_), .A2(new_n246_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n243_), .B(KEYINPUT36), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n256_), .A2(KEYINPUT37), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(KEYINPUT37), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n251_), .A2(new_n256_), .A3(KEYINPUT37), .A4(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G1gat), .B(G8gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G15gat), .B(G22gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT72), .B(G1gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G8gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n266_), .B2(KEYINPUT14), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n267_), .A2(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n263_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(KEYINPUT14), .ZN(new_n273_));
  INV_X1    g072(.A(new_n264_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT73), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n269_), .A3(new_n262_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n278_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G127gat), .B(G155gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT16), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G183gat), .B(G211gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(KEYINPUT17), .B2(new_n294_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n288_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n296_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n261_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n223_), .A2(new_n285_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n285_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n213_), .A3(new_n214_), .A4(new_n222_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(KEYINPUT12), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT12), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n223_), .A2(new_n306_), .A3(new_n285_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT64), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n304_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n310_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G120gat), .B(G148gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(G176gat), .B(G204gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n312_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT13), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n301_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT102), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G78gat), .B(G106gat), .ZN(new_n326_));
  INV_X1    g125(.A(G228gat), .ZN(new_n327_));
  INV_X1    g126(.A(G233gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT83), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(G155gat), .A3(G162gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT2), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n336_), .B1(new_n339_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT85), .B(new_n336_), .C1(new_n339_), .C2(new_n346_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n338_), .B(new_n337_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n333_), .A2(new_n335_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT1), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n331_), .B1(new_n354_), .B2(KEYINPUT1), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT84), .B1(new_n360_), .B2(new_n331_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n353_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT29), .B1(new_n351_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G197gat), .B(G204gat), .Z(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(KEYINPUT21), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(KEYINPUT21), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n330_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n334_), .B1(G155gat), .B2(G162gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n332_), .A2(KEYINPUT83), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT1), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n331_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n357_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n355_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n361_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n352_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n349_), .A2(new_n350_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n372_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n370_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n329_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n326_), .B1(new_n371_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n363_), .A2(new_n370_), .A3(new_n330_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n329_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n326_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n389_), .A3(KEYINPUT88), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n386_), .A2(new_n387_), .A3(new_n391_), .A4(new_n388_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G22gat), .B(G50gat), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n380_), .A2(new_n381_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT28), .B1(new_n396_), .B2(KEYINPUT29), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n379_), .A2(new_n352_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n372_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n398_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n395_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n401_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n400_), .B1(new_n399_), .B2(new_n372_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT86), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n394_), .A3(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n404_), .A2(KEYINPUT87), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT87), .B1(new_n404_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n393_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n389_), .B1(new_n385_), .B2(KEYINPUT89), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n386_), .A2(new_n387_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(new_n326_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n402_), .A2(new_n403_), .A3(new_n395_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n394_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G127gat), .B(G134gat), .Z(new_n428_));
  XOR2_X1   g227(.A(G113gat), .B(G120gat), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G127gat), .B(G134gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G120gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(KEYINPUT81), .A3(new_n433_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n351_), .B2(new_n362_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n380_), .A2(new_n381_), .A3(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT97), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT97), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n444_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n380_), .A2(new_n381_), .A3(new_n434_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n436_), .A2(new_n437_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT4), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n439_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n440_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n427_), .B1(new_n446_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT100), .ZN(new_n455_));
  INV_X1    g254(.A(new_n440_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n449_), .A2(KEYINPUT4), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n427_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(new_n455_), .A3(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(KEYINPUT100), .B(new_n427_), .C1(new_n446_), .C2(new_n453_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT26), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(G190gat), .ZN(new_n467_));
  INV_X1    g266(.A(G190gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT26), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT25), .B(G183gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(KEYINPUT26), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(G190gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT91), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476_));
  INV_X1    g275(.A(G169gat), .ZN(new_n477_));
  INV_X1    g276(.A(G176gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G169gat), .A2(G176gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(KEYINPUT24), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G183gat), .A2(G190gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(KEYINPUT23), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n479_), .A2(KEYINPUT24), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n476_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT93), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n475_), .A2(new_n481_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT92), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n482_), .A4(new_n489_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n497_));
  INV_X1    g296(.A(G183gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n468_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT78), .B(KEYINPUT23), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n484_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n484_), .A2(KEYINPUT23), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G169gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n478_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n480_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n497_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n510_), .B(KEYINPUT94), .C1(new_n512_), .C2(new_n500_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n492_), .A2(new_n496_), .A3(new_n514_), .A4(new_n383_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G226gat), .A2(G233gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT19), .Z(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT20), .ZN(new_n518_));
  INV_X1    g317(.A(new_n487_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n519_), .B(new_n499_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n477_), .B2(KEYINPUT22), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n478_), .B(new_n522_), .C1(new_n506_), .C2(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n523_), .A3(new_n480_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n488_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G190gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n471_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n481_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n525_), .B(new_n511_), .C1(new_n528_), .C2(KEYINPUT77), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(KEYINPUT77), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n518_), .B1(new_n531_), .B2(new_n370_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n515_), .A2(KEYINPUT95), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT95), .B1(new_n515_), .B2(new_n532_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n517_), .B(KEYINPUT90), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT20), .B1(new_n531_), .B2(new_n370_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n492_), .A2(new_n496_), .A3(new_n514_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n370_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n533_), .A2(new_n534_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT18), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G64gat), .B(G92gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  OAI221_X1 g345(.A(new_n544_), .B1(new_n539_), .B2(new_n536_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT27), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n536_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n531_), .A2(new_n370_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI22_X1  g352(.A1(new_n490_), .A2(new_n491_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT99), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n370_), .B1(new_n554_), .B2(KEYINPUT99), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n550_), .B1(new_n517_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n549_), .B1(new_n558_), .B2(new_n545_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n548_), .A2(new_n549_), .B1(new_n559_), .B2(new_n547_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n422_), .A2(new_n464_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n544_), .A2(KEYINPUT32), .ZN(new_n562_));
  OAI221_X1 g361(.A(new_n562_), .B1(new_n539_), .B2(new_n536_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n462_), .A2(new_n463_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n456_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n439_), .A2(new_n456_), .A3(new_n441_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n427_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT33), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n461_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n446_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(KEYINPUT33), .A3(new_n460_), .A4(new_n459_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n571_), .A2(new_n573_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n404_), .A2(KEYINPUT87), .A3(new_n409_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n579_), .A2(new_n393_), .B1(new_n420_), .B2(new_n417_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n561_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n438_), .B(KEYINPUT31), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G99gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT80), .B(G43gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n531_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G227gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(G15gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G71gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n588_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n588_), .B2(new_n592_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n585_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n588_), .A2(new_n592_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n596_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n588_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n584_), .A3(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n548_), .A2(new_n549_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n559_), .A2(new_n547_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(KEYINPUT101), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n555_), .A2(new_n556_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n553_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n517_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n535_), .B(new_n537_), .C1(new_n370_), .C2(new_n538_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n545_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n615_), .A2(new_n547_), .A3(KEYINPUT27), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT27), .B1(new_n546_), .B2(new_n547_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n610_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n422_), .B1(new_n609_), .B2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n605_), .A2(new_n464_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n582_), .A2(new_n606_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n272_), .A2(new_n277_), .A3(new_n229_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT75), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n272_), .A2(KEYINPUT75), .A3(new_n229_), .A4(new_n277_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n278_), .B2(new_n226_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n277_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n262_), .B1(new_n276_), .B2(new_n269_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n226_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n272_), .A2(new_n277_), .A3(new_n227_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n628_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n630_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G169gat), .B(G197gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n636_), .A3(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT76), .Z(new_n645_));
  OAI21_X1  g444(.A(new_n325_), .B1(new_n621_), .B2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n616_), .A2(new_n617_), .A3(new_n610_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n607_), .B2(new_n608_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n580_), .B(new_n620_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n412_), .A2(new_n421_), .B1(new_n463_), .B2(new_n462_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n650_), .A2(new_n560_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n651_), .B2(new_n605_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n645_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT102), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n324_), .B1(new_n646_), .B2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n464_), .A2(new_n265_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT38), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT38), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n255_), .B(KEYINPUT103), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n621_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n323_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n644_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n663_), .A2(new_n300_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n666_), .B2(new_n464_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n658_), .A2(new_n659_), .A3(new_n667_), .ZN(G1324gat));
  INV_X1    g467(.A(G8gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n647_), .A2(new_n648_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n655_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  INV_X1    g471(.A(new_n666_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(KEYINPUT104), .A3(new_n670_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  INV_X1    g474(.A(new_n670_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n666_), .B2(new_n676_), .ZN(new_n677_));
  AND4_X1   g476(.A1(new_n672_), .A2(new_n674_), .A3(G8gat), .A4(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n666_), .A2(new_n676_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n669_), .B1(new_n679_), .B2(KEYINPUT104), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n672_), .B1(new_n680_), .B2(new_n677_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n671_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT40), .B(new_n671_), .C1(new_n678_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1325gat));
  OAI21_X1  g485(.A(G15gat), .B1(new_n666_), .B2(new_n606_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT41), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n655_), .A2(new_n594_), .A3(new_n605_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n666_), .B2(new_n580_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT42), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n580_), .A2(G22gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT105), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n655_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n299_), .A2(new_n255_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n323_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n646_), .B2(new_n654_), .ZN(new_n699_));
  INV_X1    g498(.A(G29gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n464_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n699_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n323_), .A2(new_n644_), .A3(new_n300_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n261_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n621_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n652_), .A2(new_n706_), .A3(new_n261_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n464_), .B1(new_n708_), .B2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT107), .B1(new_n714_), .B2(G29gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n716_), .B(new_n700_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n702_), .B1(new_n715_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n646_), .A2(new_n654_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n698_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n676_), .A2(G36gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n699_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(KEYINPUT45), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n708_), .A2(KEYINPUT44), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n670_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n712_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n719_), .B1(new_n731_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n711_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n710_), .B1(new_n708_), .B2(KEYINPUT106), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G36gat), .B1(new_n740_), .B2(new_n734_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT46), .A3(new_n730_), .A4(new_n729_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1329gat));
  INV_X1    g542(.A(G43gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n606_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n712_), .A2(new_n733_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n699_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n747_), .B2(new_n606_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(KEYINPUT47), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT47), .B1(new_n746_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n699_), .B2(new_n422_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n733_), .A2(G50gat), .A3(new_n422_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n712_), .B2(new_n753_), .ZN(G1331gat));
  NOR3_X1   g553(.A1(new_n653_), .A2(new_n323_), .A3(new_n300_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n662_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n464_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n652_), .A2(new_n664_), .A3(new_n663_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n300_), .A3(new_n261_), .ZN(new_n760_));
  INV_X1    g559(.A(G57gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n701_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n756_), .B2(new_n670_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT48), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n764_), .A3(new_n670_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n756_), .B2(new_n605_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n760_), .A2(new_n769_), .A3(new_n605_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n756_), .B2(new_n422_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT50), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n760_), .A2(new_n775_), .A3(new_n422_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1335gat));
  NOR3_X1   g578(.A1(new_n323_), .A2(new_n299_), .A3(new_n644_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n464_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n759_), .A2(new_n299_), .A3(new_n255_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n215_), .A3(new_n701_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT110), .ZN(G1336gat));
  OAI21_X1  g587(.A(G92gat), .B1(new_n783_), .B2(new_n676_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n216_), .A3(new_n670_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n783_), .B2(new_n606_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(new_n605_), .A3(new_n219_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n785_), .A2(new_n206_), .A3(new_n422_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n580_), .B(new_n781_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n206_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n652_), .A2(new_n706_), .A3(new_n261_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n706_), .B1(new_n652_), .B2(new_n261_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n422_), .B(new_n780_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT111), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n797_), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G106gat), .B1(new_n803_), .B2(KEYINPUT111), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n782_), .B2(new_n422_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(KEYINPUT52), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n796_), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n796_), .C1(new_n805_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n312_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n310_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT55), .B1(new_n817_), .B2(KEYINPUT113), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n816_), .B(new_n818_), .C1(new_n311_), .C2(new_n308_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n319_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n312_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n626_), .A2(new_n633_), .A3(new_n628_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n640_), .B1(new_n635_), .B2(new_n627_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n643_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n823_), .A2(new_n643_), .A3(new_n826_), .A4(KEYINPUT116), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n308_), .A2(new_n311_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n308_), .B2(new_n311_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n815_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n319_), .B1(new_n834_), .B2(new_n818_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n831_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n261_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n829_), .A2(new_n830_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n840_), .B2(new_n822_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n320_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(KEYINPUT114), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n835_), .B2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n319_), .B(new_n844_), .C1(new_n834_), .C2(new_n818_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT115), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n821_), .A2(new_n844_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n835_), .A2(new_n845_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .A4(new_n843_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n322_), .A2(new_n643_), .A3(new_n826_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n255_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n842_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(KEYINPUT57), .A3(new_n255_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n299_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n324_), .B2(new_n653_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n301_), .A2(new_n645_), .A3(new_n323_), .A4(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT117), .B1(new_n859_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n861_), .A2(new_n864_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n854_), .A2(KEYINPUT57), .A3(new_n255_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n854_), .B2(new_n255_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n842_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n867_), .B(new_n868_), .C1(new_n871_), .C2(new_n299_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n619_), .A2(new_n701_), .A3(new_n605_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n876_), .B(new_n299_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n855_), .A2(new_n856_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n842_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n858_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n880_), .B2(new_n300_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n868_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n873_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n873_), .A2(new_n883_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n875_), .A2(new_n653_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G113gat), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n874_), .A2(G113gat), .A3(new_n664_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1340gat));
  NAND3_X1  g691(.A1(new_n875_), .A2(new_n663_), .A3(new_n888_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G120gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895_));
  AOI21_X1  g694(.A(G120gat), .B1(new_n663_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n895_), .B2(G120gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI211_X1 g697(.A(KEYINPUT121), .B(G120gat), .C1(new_n663_), .C2(new_n895_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n874_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n900_), .ZN(G1341gat));
  NAND3_X1  g700(.A1(new_n875_), .A2(new_n299_), .A3(new_n888_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G127gat), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n874_), .A2(G127gat), .A3(new_n300_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1342gat));
  INV_X1    g704(.A(G134gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n874_), .B2(new_n660_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT122), .B(new_n906_), .C1(new_n874_), .C2(new_n660_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n874_), .A2(KEYINPUT59), .B1(new_n882_), .B2(new_n887_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n704_), .A2(new_n906_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1343gat));
  AND2_X1   g712(.A1(new_n866_), .A2(new_n872_), .ZN(new_n914_));
  NOR4_X1   g713(.A1(new_n670_), .A2(new_n464_), .A3(new_n580_), .A4(new_n605_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n644_), .A3(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n663_), .A3(new_n915_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g718(.A1(new_n914_), .A2(new_n299_), .A3(new_n915_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  INV_X1    g721(.A(G162gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n914_), .A2(new_n923_), .A3(new_n661_), .A4(new_n915_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n914_), .A2(new_n261_), .A3(new_n915_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1347gat));
  INV_X1    g725(.A(new_n882_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n670_), .A2(new_n620_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n422_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n927_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n644_), .A2(new_n506_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT124), .Z(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n882_), .A2(new_n644_), .A3(new_n929_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n936_));
  AND3_X1   g735(.A1(new_n935_), .A2(G169gat), .A3(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n935_), .B2(G169gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n934_), .B1(new_n937_), .B2(new_n938_), .ZN(G1348gat));
  AND2_X1   g738(.A1(new_n914_), .A2(new_n580_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n928_), .A2(new_n478_), .A3(new_n323_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n882_), .A2(new_n663_), .A3(new_n929_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n940_), .A2(new_n941_), .B1(new_n942_), .B2(new_n478_), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n300_), .A2(new_n471_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n928_), .A2(new_n300_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n914_), .A2(new_n580_), .A3(new_n945_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n931_), .A2(new_n944_), .B1(new_n946_), .B2(new_n498_), .ZN(G1350gat));
  AND2_X1   g746(.A1(new_n470_), .A2(new_n474_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n931_), .A2(new_n948_), .A3(new_n661_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n927_), .A2(new_n704_), .A3(new_n930_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n468_), .B2(new_n950_), .ZN(G1351gat));
  AND3_X1   g750(.A1(new_n670_), .A2(new_n650_), .A3(new_n606_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n866_), .A2(new_n644_), .A3(new_n872_), .A4(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(G197gat), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(KEYINPUT126), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n953_), .A2(new_n957_), .A3(new_n954_), .ZN(new_n958_));
  AND3_X1   g757(.A1(new_n866_), .A2(new_n872_), .A3(new_n952_), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n959_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n644_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n962_));
  AOI22_X1  g761(.A1(new_n956_), .A2(new_n958_), .B1(new_n960_), .B2(new_n962_), .ZN(G1352gat));
  NAND2_X1  g762(.A1(new_n959_), .A2(new_n663_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT127), .B(G204gat), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n964_), .B(new_n965_), .ZN(G1353gat));
  OR2_X1    g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n959_), .B2(new_n299_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n959_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n300_), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT63), .B(G211gat), .Z(new_n971_));
  AOI21_X1  g770(.A(new_n968_), .B1(new_n970_), .B2(new_n971_), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n969_), .B2(new_n704_), .ZN(new_n973_));
  OR2_X1    g772(.A1(new_n660_), .A2(G218gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n969_), .B2(new_n974_), .ZN(G1355gat));
endmodule


