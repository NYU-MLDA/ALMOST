//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n212_), .A2(KEYINPUT77), .A3(KEYINPUT22), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT78), .B(G176gat), .Z(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT22), .B1(new_n212_), .B2(KEYINPUT77), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n210_), .B(new_n211_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n220_), .A2(new_n209_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT22), .B(G169gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n214_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n224_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n226_), .B(KEYINPUT20), .C1(new_n207_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G226gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT19), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n207_), .A2(new_n231_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(KEYINPUT20), .C1(new_n207_), .C2(new_n225_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n240_));
  XNOR2_X1  g039(.A(G8gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G64gat), .B(G92gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n235_), .A2(new_n246_), .A3(new_n238_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n232_), .A2(new_n234_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT96), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n249_), .B1(new_n247_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n256_), .B2(new_n247_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n250_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G155gat), .B(G162gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT81), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  OAI22_X1  g067(.A1(new_n263_), .A2(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n267_), .B(KEYINPUT79), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT82), .B(KEYINPUT2), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n262_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(KEYINPUT1), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n277_), .A2(KEYINPUT80), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n275_), .A2(KEYINPUT1), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n277_), .B2(KEYINPUT80), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n274_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n273_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT84), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n285_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n273_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT91), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT90), .B(KEYINPUT4), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n288_), .A4(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n283_), .A2(new_n285_), .A3(new_n288_), .A4(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT91), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n302_), .B(new_n304_), .C1(new_n305_), .C2(new_n292_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n296_), .B1(new_n306_), .B2(new_n295_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT94), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT93), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n316_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n309_), .B1(new_n307_), .B2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n259_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n283_), .A2(new_n285_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AOI211_X1 g125(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n283_), .C2(new_n285_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT85), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT28), .B1(new_n299_), .B2(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  AND3_X1   g132(.A1(new_n328_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n322_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(new_n332_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT88), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(G233gat), .ZN(new_n343_));
  OAI221_X1 g142(.A(new_n207_), .B1(new_n342_), .B2(new_n343_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT29), .B1(new_n273_), .B2(new_n281_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n207_), .A3(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n342_), .A2(new_n343_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n349_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n207_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n345_), .B(new_n351_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n344_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n344_), .C1(new_n352_), .C2(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n336_), .A2(new_n341_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n339_), .A2(new_n340_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n364_), .A2(new_n322_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n225_), .B(KEYINPUT30), .ZN(new_n366_));
  XOR2_X1   g165(.A(G71gat), .B(G99gat), .Z(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n366_), .B(new_n369_), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n290_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT31), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n366_), .B(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n288_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n371_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n373_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n363_), .A2(new_n365_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n321_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n246_), .A2(KEYINPUT32), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n239_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n382_), .B2(new_n252_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n320_), .A2(new_n317_), .A3(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n306_), .A2(new_n295_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n316_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n248_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT33), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n307_), .A2(KEYINPUT33), .A3(new_n315_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n378_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n381_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G8gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G1gat), .ZN(new_n401_));
  INV_X1    g200(.A(G8gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT14), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G22gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n403_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G29gat), .B(G36gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G43gat), .B(G50gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G29gat), .B(G36gat), .Z(new_n412_));
  XOR2_X1   g211(.A(G43gat), .B(G50gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n411_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(G229gat), .A3(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT15), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(KEYINPUT15), .A3(new_n411_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n408_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G229gat), .A2(G233gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT74), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n417_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G113gat), .B(G141gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G169gat), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n419_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT75), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n419_), .A2(new_n434_), .A3(new_n427_), .A4(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(new_n427_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(KEYINPUT76), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(KEYINPUT76), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n398_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G230gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(new_n343_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G85gat), .B(G92gat), .Z(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n453_), .B2(KEYINPUT9), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n454_), .B(new_n457_), .C1(KEYINPUT9), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT8), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT64), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n450_), .A2(new_n451_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n456_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT64), .A3(new_n462_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n460_), .B1(new_n471_), .B2(new_n453_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n462_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n452_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n453_), .A2(new_n460_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n459_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(KEYINPUT11), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT65), .B(new_n459_), .C1(new_n472_), .C2(new_n476_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n479_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n447_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G120gat), .B(G148gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G204gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT5), .B(G176gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND3_X1  g292(.A1(new_n479_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n484_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n494_), .B(new_n495_), .C1(new_n488_), .C2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n489_), .B(new_n493_), .C1(new_n498_), .C2(new_n447_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n494_), .A2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n453_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n452_), .B1(new_n473_), .B2(new_n461_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(new_n470_), .ZN(new_n505_));
  OAI22_X1  g304(.A1(new_n505_), .A2(new_n460_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT65), .B1(new_n506_), .B2(new_n459_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n486_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n484_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n447_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n512_), .A2(KEYINPUT67), .A3(new_n489_), .A4(new_n493_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n501_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n489_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n493_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT68), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT13), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n514_), .A2(new_n517_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G127gat), .B(G155gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT16), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G183gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n525_), .B(KEYINPUT16), .ZN(new_n528_));
  INV_X1    g327(.A(G183gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n530_), .A3(G211gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(G211gat), .B1(new_n527_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT17), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n408_), .A2(KEYINPUT72), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n538_));
  INV_X1    g337(.A(G231gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(new_n343_), .ZN(new_n540_));
  OR3_X1    g339(.A1(new_n536_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n540_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n541_), .A2(new_n484_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n484_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n532_), .A2(KEYINPUT17), .A3(new_n533_), .ZN(new_n545_));
  NOR4_X1   g344(.A1(new_n535_), .A2(new_n543_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n535_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n535_), .B(KEYINPUT73), .C1(new_n543_), .C2(new_n544_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n479_), .A2(new_n416_), .A3(new_n486_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n421_), .A2(new_n422_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n477_), .A2(new_n555_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(new_n556_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n554_), .B(new_n560_), .C1(new_n556_), .C2(new_n559_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G190gat), .B(G218gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT69), .Z(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT70), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n563_), .A2(new_n573_), .A3(new_n564_), .A4(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n563_), .A2(new_n564_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n567_), .B(KEYINPUT36), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT71), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n553_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n577_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n582_));
  AOI211_X1 g381(.A(KEYINPUT37), .B(new_n582_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n524_), .A2(new_n552_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n445_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n320_), .A2(new_n317_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n401_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n440_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n524_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n551_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n582_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n398_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n597_), .B2(new_n587_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n589_), .A2(new_n590_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n591_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT97), .ZN(G1324gat));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n259_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(G8gat), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(new_n259_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(G8gat), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n604_), .A2(new_n605_), .B1(new_n586_), .B2(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n604_), .A2(new_n605_), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT98), .B(new_n402_), .C1(new_n596_), .C2(new_n259_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n596_), .B2(new_n394_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n586_), .A2(new_n614_), .A3(new_n394_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n363_), .A2(new_n365_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n596_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n586_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(G29gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n593_), .A2(new_n552_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n397_), .B2(new_n584_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n584_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT43), .B(new_n631_), .C1(new_n381_), .C2(new_n396_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT44), .B(new_n628_), .C1(new_n630_), .C2(new_n632_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n588_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n626_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n638_), .B2(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n552_), .A2(new_n595_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n524_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n445_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n587_), .A2(G29gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT101), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n640_), .B1(new_n643_), .B2(new_n645_), .ZN(G1328gat));
  NOR2_X1   g445(.A1(new_n606_), .A2(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n445_), .A2(new_n642_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n635_), .A2(new_n259_), .A3(new_n636_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G36gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT46), .B(new_n649_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  AND2_X1   g457(.A1(new_n394_), .A2(G43gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n635_), .A2(new_n636_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n635_), .A2(new_n662_), .A3(new_n636_), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(G43gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n643_), .B2(new_n378_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT47), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n669_), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1330gat));
  NAND4_X1  g470(.A1(new_n635_), .A2(G50gat), .A3(new_n621_), .A4(new_n636_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n643_), .A2(new_n620_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(G50gat), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT105), .Z(G1331gat));
  INV_X1    g474(.A(G57gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n523_), .A2(new_n440_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n397_), .A2(new_n551_), .A3(new_n631_), .A4(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n678_), .B2(new_n587_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT106), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n398_), .A2(new_n595_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n551_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n523_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n684_), .A2(new_n676_), .A3(new_n587_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n680_), .A2(new_n685_), .ZN(G1332gat));
  OR3_X1    g485(.A1(new_n678_), .A2(G64gat), .A3(new_n606_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G64gat), .B1(new_n684_), .B2(new_n606_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT107), .ZN(G1333gat));
  OAI21_X1  g491(.A(G71gat), .B1(new_n684_), .B2(new_n378_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT49), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n378_), .A2(G71gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n678_), .B2(new_n695_), .ZN(G1334gat));
  OAI21_X1  g495(.A(G78gat), .B1(new_n684_), .B2(new_n620_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT50), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n620_), .A2(G78gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n678_), .B2(new_n699_), .ZN(G1335gat));
  INV_X1    g499(.A(new_n677_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n551_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n587_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n398_), .A2(new_n641_), .A3(new_n701_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n587_), .A2(G85gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(G92gat), .B1(new_n703_), .B2(new_n606_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n606_), .A2(G92gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n706_), .B2(new_n710_), .ZN(G1337gat));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n394_), .A3(new_n455_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n703_), .A2(new_n378_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G99gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G99gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g517(.A1(new_n705_), .A2(new_n456_), .A3(new_n621_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n703_), .A2(new_n620_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G106gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G106gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g524(.A(G113gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT59), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n592_), .B1(new_n501_), .B2(new_n513_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n498_), .B2(new_n447_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n511_), .A2(KEYINPUT110), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n498_), .B2(new_n731_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n733_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n502_), .A2(new_n510_), .A3(KEYINPUT55), .A4(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n516_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n730_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n418_), .A2(new_n426_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n423_), .A2(new_n417_), .A3(new_n425_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n438_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n436_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n744_), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT111), .B(new_n746_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n595_), .B1(new_n740_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n729_), .B1(new_n751_), .B2(KEYINPUT57), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n737_), .A2(new_n516_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n749_), .B1(new_n758_), .B2(new_n730_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT112), .B(new_n753_), .C1(new_n759_), .C2(new_n595_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n748_), .B1(new_n501_), .B2(new_n513_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(KEYINPUT58), .C1(new_n738_), .C2(new_n739_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n745_), .A2(new_n747_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n514_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT113), .B(KEYINPUT58), .Z(new_n766_));
  OAI211_X1 g565(.A(new_n584_), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n751_), .A2(KEYINPUT57), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n752_), .A2(new_n760_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n552_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n682_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n551_), .A2(new_n441_), .A3(KEYINPUT109), .A4(new_n442_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n584_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n523_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(new_n523_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n770_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n588_), .A2(new_n606_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n380_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n728_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n728_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n767_), .B(KEYINPUT114), .C1(KEYINPUT57), .C2(new_n751_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n768_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n753_), .B1(new_n759_), .B2(new_n595_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT114), .B1(new_n790_), .B2(new_n767_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n552_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n787_), .B1(new_n792_), .B2(new_n780_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n727_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n779_), .B1(new_n769_), .B2(new_n552_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n784_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  INV_X1    g596(.A(new_n767_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n740_), .A2(new_n750_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n595_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n768_), .A3(new_n788_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n779_), .B1(new_n803_), .B2(new_n552_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n796_), .B(KEYINPUT115), .C1(new_n804_), .C2(new_n787_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n794_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n726_), .B1(new_n806_), .B2(new_n443_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n781_), .A2(new_n785_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n440_), .A2(new_n726_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT116), .B1(new_n807_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n444_), .B1(new_n794_), .B2(new_n805_), .ZN(new_n813_));
  OAI221_X1 g612(.A(new_n812_), .B1(new_n808_), .B2(new_n809_), .C1(new_n813_), .C2(new_n726_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(G1340gat));
  NOR2_X1   g614(.A1(new_n795_), .A2(new_n784_), .ZN(new_n816_));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n523_), .B2(KEYINPUT60), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n816_), .B(new_n818_), .C1(KEYINPUT60), .C2(new_n817_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT117), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n786_), .A2(new_n793_), .A3(new_n523_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n817_), .B2(new_n821_), .ZN(G1341gat));
  INV_X1    g621(.A(new_n806_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G127gat), .B1(new_n823_), .B2(new_n552_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n552_), .A2(G127gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n808_), .B2(new_n825_), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n823_), .B2(new_n631_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n800_), .A2(G134gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n808_), .B2(new_n828_), .ZN(G1343gat));
  INV_X1    g628(.A(new_n379_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n795_), .A2(new_n830_), .A3(new_n782_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n440_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT118), .B(G141gat), .Z(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1344gat));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n524_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT119), .B(G148gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1345gat));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n838_), .A3(new_n551_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n831_), .B2(new_n551_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT61), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n839_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n842_), .A2(new_n845_), .A3(G155gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(G155gat), .B1(new_n842_), .B2(new_n845_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n795_), .A2(new_n830_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n783_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n851_), .B2(new_n800_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT121), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n851_), .A2(new_n849_), .A3(new_n631_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1347gat));
  NOR3_X1   g654(.A1(new_n588_), .A2(new_n378_), .A3(new_n606_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n620_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n804_), .A2(KEYINPUT123), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT123), .B1(new_n804_), .B2(new_n857_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n858_), .A2(new_n228_), .A3(new_n440_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n792_), .A2(new_n780_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n857_), .A2(new_n592_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n212_), .B1(new_n864_), .B2(KEYINPUT122), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n866_), .A3(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n861_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n863_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT122), .B1(new_n804_), .B2(new_n869_), .ZN(new_n870_));
  AND4_X1   g669(.A1(new_n861_), .A2(new_n870_), .A3(new_n867_), .A4(G169gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n860_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n860_), .C1(new_n868_), .C2(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n781_), .A2(new_n620_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n856_), .A2(G176gat), .A3(new_n524_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n858_), .A2(new_n524_), .A3(new_n859_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n214_), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n856_), .A2(new_n551_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n529_), .B1(new_n877_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n858_), .A2(new_n859_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n552_), .A2(new_n218_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n884_), .B2(new_n631_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n595_), .A2(new_n219_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n884_), .B2(new_n890_), .ZN(G1351gat));
  NOR2_X1   g690(.A1(new_n588_), .A2(new_n606_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n850_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n440_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n430_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n895_), .A2(new_n430_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(G1352gat));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n524_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g701(.A(new_n552_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(new_n904_));
  NAND2_X1  g703(.A1(new_n894_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n905_), .B(new_n906_), .Z(G1354gat));
  OR3_X1    g706(.A1(new_n893_), .A2(G218gat), .A3(new_n800_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G218gat), .B1(new_n893_), .B2(new_n631_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1355gat));
endmodule


