//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G85gat), .A3(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G85gat), .B(G92gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n204_), .B(new_n206_), .C1(new_n205_), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT10), .B(G99gat), .Z(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT65), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  AOI211_X1 g016(.A(KEYINPUT8), .B(new_n207_), .C1(new_n217_), .C2(new_n204_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n207_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n204_), .A2(KEYINPUT66), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n217_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n204_), .A2(KEYINPUT66), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n218_), .B1(new_n223_), .B2(KEYINPUT8), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n213_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT72), .B(G43gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G50gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G232gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT71), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT34), .ZN(new_n235_));
  INV_X1    g034(.A(new_n230_), .ZN(new_n236_));
  OAI221_X1 g035(.A(new_n232_), .B1(KEYINPUT35), .B2(new_n235_), .C1(new_n226_), .C2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(KEYINPUT35), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT36), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G190gat), .B(G218gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G134gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(G162gat), .Z(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n242_), .B1(new_n241_), .B2(new_n245_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n202_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(KEYINPUT37), .A3(new_n248_), .A4(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT74), .B(G8gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G1gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT14), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G15gat), .B(G22gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT75), .ZN(new_n260_));
  INV_X1    g059(.A(G1gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G8gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT67), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT11), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G71gat), .B(G78gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n266_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n264_), .B(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G127gat), .B(G155gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G183gat), .B(G211gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT17), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n281_), .B(KEYINPUT17), .Z(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n276_), .B2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n254_), .A2(KEYINPUT77), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT77), .B1(new_n254_), .B2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n225_), .A2(new_n273_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT12), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n272_), .B(new_n270_), .C1(new_n213_), .C2(new_n224_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  AND2_X1   g090(.A1(G230gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(KEYINPUT68), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G120gat), .B(G148gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G176gat), .B(G204gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT70), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n294_), .A2(new_n303_), .A3(new_n297_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT13), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT13), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n286_), .A2(new_n287_), .A3(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT78), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT3), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT2), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n316_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(KEYINPUT1), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n318_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G22gat), .B(G50gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT28), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n331_), .B(new_n333_), .Z(new_n334_));
  XOR2_X1   g133(.A(G78gat), .B(G106gat), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n331_), .B(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(KEYINPUT88), .B2(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT86), .B1(new_n342_), .B2(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(KEYINPUT21), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n347_));
  XOR2_X1   g146(.A(G197gat), .B(G204gat), .Z(new_n348_));
  NAND4_X1  g147(.A1(new_n348_), .A2(KEYINPUT21), .A3(new_n341_), .A4(new_n343_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G233gat), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n352_), .A2(KEYINPUT85), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(KEYINPUT85), .ZN(new_n354_));
  OAI21_X1  g153(.A(G228gat), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n351_), .B(new_n355_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n329_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n359_), .B2(new_n355_), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n340_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364_));
  INV_X1    g163(.A(G113gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G120gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT95), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT96), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n367_), .B(new_n329_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n368_), .B(new_n371_), .C1(new_n373_), .C2(new_n363_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G85gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT33), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT18), .B(G64gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G169gat), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(G190gat), .ZN(new_n395_));
  INV_X1    g194(.A(G183gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G190gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT23), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n394_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n412_), .B2(KEYINPUT26), .ZN(new_n413_));
  NAND2_X1  g212(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT25), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n408_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n390_), .A2(KEYINPUT24), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT82), .B1(new_n417_), .B2(new_n406_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT24), .A4(new_n390_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n402_), .A2(KEYINPUT83), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(new_n401_), .A3(G183gat), .A4(G190gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n400_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n405_), .B1(new_n416_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n389_), .B1(new_n428_), .B2(new_n351_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT25), .B(G183gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n432_), .A2(new_n409_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT26), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n399_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT90), .B1(new_n436_), .B2(new_n431_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n430_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n419_), .A3(new_n390_), .A4(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n419_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n403_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n396_), .A2(new_n399_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n426_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n446_), .A2(KEYINPUT92), .A3(new_n394_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT92), .B1(new_n446_), .B2(new_n394_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n350_), .B(new_n444_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(KEYINPUT89), .Z(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT19), .Z(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n429_), .A2(new_n449_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n429_), .A2(new_n449_), .A3(KEYINPUT93), .A4(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n389_), .B1(new_n459_), .B2(new_n351_), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n393_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n390_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n403_), .B2(new_n397_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n422_), .A2(new_n426_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n436_), .B1(new_n395_), .B2(new_n435_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n414_), .B(KEYINPUT25), .Z(new_n468_));
  AOI22_X1  g267(.A1(new_n467_), .A2(new_n468_), .B1(new_n407_), .B2(new_n406_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n350_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n453_), .B1(new_n460_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n388_), .B1(new_n458_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n446_), .A2(new_n394_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n446_), .A2(KEYINPUT92), .A3(new_n394_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n438_), .A2(new_n403_), .A3(new_n443_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n476_), .A2(new_n477_), .B1(new_n478_), .B2(new_n441_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT20), .B(new_n471_), .C1(new_n479_), .C2(new_n350_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n452_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n481_), .A2(new_n387_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(KEYINPUT94), .A3(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n458_), .A2(new_n472_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT94), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n387_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n381_), .B1(new_n372_), .B2(new_n371_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n368_), .B1(new_n373_), .B2(new_n363_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n370_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n383_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n374_), .A2(new_n376_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n380_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n382_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n460_), .A2(new_n453_), .A3(new_n471_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n444_), .A2(new_n350_), .A3(new_n474_), .ZN(new_n497_));
  AOI211_X1 g296(.A(new_n496_), .B(new_n453_), .C1(new_n429_), .C2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n497_), .B(KEYINPUT20), .C1(new_n470_), .C2(new_n350_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT97), .B1(new_n499_), .B2(new_n452_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n495_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT32), .A3(new_n387_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n484_), .B1(new_n503_), .B2(new_n388_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n362_), .B1(new_n491_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n483_), .A2(new_n507_), .A3(new_n486_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n501_), .A2(KEYINPUT98), .A3(new_n388_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT98), .B1(new_n501_), .B2(new_n388_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT27), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n482_), .B(KEYINPUT99), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT100), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n501_), .A2(new_n388_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n501_), .A2(KEYINPUT98), .A3(new_n388_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n458_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n519_), .A2(KEYINPUT99), .A3(new_n387_), .A4(new_n481_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT99), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n482_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT100), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n518_), .A2(new_n523_), .A3(new_n524_), .A4(KEYINPUT27), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n508_), .B(new_n361_), .C1(new_n513_), .C2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n494_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n506_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n428_), .B(KEYINPUT30), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT84), .ZN(new_n530_));
  XOR2_X1   g329(.A(G15gat), .B(G43gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G227gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT31), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n367_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n529_), .A2(KEYINPUT84), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT101), .B1(new_n528_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n513_), .A2(new_n525_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n508_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n362_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n527_), .A3(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n543_), .A2(new_n527_), .A3(new_n544_), .A4(new_n362_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n491_), .A2(new_n505_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n362_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT101), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n540_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n262_), .B(G8gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n230_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n264_), .A2(new_n231_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n264_), .A2(new_n236_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G169gat), .B(G197gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G141gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT79), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n365_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n558_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n314_), .B2(KEYINPUT78), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n315_), .A2(new_n553_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n261_), .A3(new_n494_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT104), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n572_), .A2(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(KEYINPUT104), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT103), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n252_), .A2(KEYINPUT103), .A3(new_n248_), .A4(new_n246_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n285_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n553_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n585_), .A2(new_n313_), .A3(new_n569_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G1gat), .B1(new_n587_), .B2(new_n527_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .A4(new_n588_), .ZN(G1324gat));
  INV_X1    g388(.A(new_n545_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n255_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n571_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G8gat), .B1(new_n587_), .B2(new_n590_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g396(.A(KEYINPUT105), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n586_), .A2(new_n541_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(G15gat), .ZN(new_n600_));
  INV_X1    g399(.A(G15gat), .ZN(new_n601_));
  AOI211_X1 g400(.A(KEYINPUT105), .B(new_n601_), .C1(new_n586_), .C2(new_n541_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT41), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n571_), .A2(new_n601_), .A3(new_n541_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT106), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(G22gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n586_), .B2(new_n362_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT42), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n571_), .A2(new_n610_), .A3(new_n362_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1327gat));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n251_), .A2(new_n253_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n553_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT108), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n553_), .A2(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT43), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT108), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n553_), .A2(new_n621_), .A3(new_n616_), .A4(new_n615_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n312_), .A2(new_n583_), .A3(new_n568_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT107), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(KEYINPUT44), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n494_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT44), .B1(new_n623_), .B2(new_n625_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G29gat), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n553_), .A2(new_n582_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n527_), .A2(G29gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT109), .Z(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n632_), .B2(new_n634_), .ZN(G1328gat));
  NOR3_X1   g434(.A1(new_n632_), .A2(G36gat), .A3(new_n590_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT45), .Z(new_n637_));
  NAND2_X1  g436(.A1(new_n626_), .A2(new_n545_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G36gat), .B1(new_n638_), .B2(new_n628_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT110), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1329gat));
  INV_X1    g441(.A(KEYINPUT47), .ZN(new_n643_));
  INV_X1    g442(.A(new_n632_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G43gat), .B1(new_n644_), .B2(new_n541_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n626_), .A2(G43gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n623_), .A2(new_n625_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n540_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT111), .B(new_n645_), .C1(new_n646_), .C2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT111), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n648_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n652_), .A2(G43gat), .A3(new_n541_), .A4(new_n626_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n645_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n643_), .B1(new_n650_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n626_), .A2(G43gat), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n657_), .A2(new_n540_), .A3(new_n628_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT111), .B1(new_n658_), .B2(new_n645_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(KEYINPUT47), .A3(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n656_), .A2(new_n661_), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n644_), .B2(new_n362_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n626_), .A2(G50gat), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n628_), .A2(new_n361_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(G1331gat));
  NOR2_X1   g465(.A1(new_n286_), .A2(new_n287_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n312_), .A2(new_n568_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n553_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G57gat), .B1(new_n670_), .B2(new_n494_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n668_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT112), .B1(new_n585_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT112), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n584_), .A2(new_n553_), .A3(new_n674_), .A4(new_n668_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n527_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n671_), .B1(new_n677_), .B2(G57gat), .ZN(G1332gat));
  OR3_X1    g477(.A1(new_n669_), .A2(G64gat), .A3(new_n590_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G64gat), .B1(new_n676_), .B2(new_n590_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(KEYINPUT113), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(KEYINPUT113), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT48), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT48), .B1(new_n681_), .B2(new_n682_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n683_), .B2(new_n684_), .ZN(G1333gat));
  OR3_X1    g484(.A1(new_n669_), .A2(G71gat), .A3(new_n540_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G71gat), .B1(new_n676_), .B2(new_n540_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT49), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT49), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1334gat));
  OR3_X1    g489(.A1(new_n669_), .A2(G78gat), .A3(new_n361_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G78gat), .B1(new_n676_), .B2(new_n361_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT50), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT50), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(G1335gat));
  NOR2_X1   g494(.A1(new_n672_), .A2(new_n285_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n630_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n494_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n623_), .A2(new_n696_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(KEYINPUT114), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n623_), .B2(new_n696_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n527_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n698_), .B1(new_n704_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g504(.A(G92gat), .B1(new_n697_), .B2(new_n545_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n703_), .A2(new_n590_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g507(.A(KEYINPUT117), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n697_), .A2(new_n210_), .A3(new_n541_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT115), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n700_), .A2(new_n540_), .A3(new_n702_), .ZN(new_n712_));
  INV_X1    g511(.A(G99gat), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n709_), .B(new_n711_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT116), .ZN(new_n715_));
  NAND2_X1  g514(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n711_), .B(new_n716_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n715_), .A2(new_n717_), .B1(new_n718_), .B2(new_n714_), .ZN(G1338gat));
  OAI21_X1  g518(.A(G106gat), .B1(new_n699_), .B2(new_n361_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT118), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT118), .B(G106gat), .C1(new_n699_), .C2(new_n361_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT52), .A3(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n697_), .A2(new_n209_), .A3(new_n362_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n721_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n725_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n724_), .A2(new_n730_), .A3(new_n725_), .A4(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  NAND3_X1  g531(.A1(new_n285_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n309_), .A2(new_n311_), .B1(KEYINPUT119), .B2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(KEYINPUT119), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(KEYINPUT120), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT120), .B1(new_n734_), .B2(new_n735_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n254_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT54), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT54), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n582_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n568_), .A2(new_n307_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n291_), .A2(new_n744_), .A3(new_n293_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n746_));
  OAI22_X1  g545(.A1(new_n745_), .A2(new_n746_), .B1(new_n293_), .B2(new_n291_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n305_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n743_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n555_), .A2(new_n559_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n557_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n555_), .A2(new_n556_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n754_), .B(new_n565_), .C1(new_n557_), .C2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n566_), .A2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n308_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n742_), .B(KEYINPUT57), .C1(new_n752_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n752_), .A2(new_n758_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n582_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n751_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n747_), .B2(new_n305_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n307_), .B(new_n757_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n751_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(KEYINPUT58), .A3(new_n307_), .A4(new_n757_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n769_), .A3(new_n616_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n759_), .A2(new_n762_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n583_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n741_), .A2(new_n772_), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n540_), .A2(new_n545_), .A3(new_n527_), .A4(new_n362_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT59), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n771_), .A2(KEYINPUT121), .A3(new_n583_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT121), .B1(new_n771_), .B2(new_n583_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n741_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n774_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n782_));
  OAI21_X1  g581(.A(G113gat), .B1(new_n569_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n365_), .A2(KEYINPUT122), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n776_), .A2(new_n781_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n365_), .B1(new_n775_), .B2(new_n569_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1340gat));
  NAND2_X1  g586(.A1(new_n776_), .A2(new_n781_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G120gat), .B1(new_n788_), .B2(new_n312_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n775_), .ZN(new_n790_));
  INV_X1    g589(.A(G120gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n312_), .B2(KEYINPUT60), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n792_), .C1(KEYINPUT60), .C2(new_n791_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(G127gat), .B1(new_n790_), .B2(new_n285_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n776_), .A2(new_n781_), .A3(G127gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n285_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n790_), .B2(new_n582_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n776_), .A2(new_n781_), .A3(G134gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n616_), .ZN(G1343gat));
  AOI21_X1  g599(.A(new_n541_), .B1(new_n741_), .B2(new_n772_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n545_), .A2(new_n527_), .A3(new_n361_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n568_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n313_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n285_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT61), .B(G155gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  NAND4_X1  g609(.A1(new_n801_), .A2(G162gat), .A3(new_n616_), .A4(new_n802_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n801_), .A2(new_n582_), .A3(new_n802_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G162gat), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n811_), .B(KEYINPUT123), .C1(new_n812_), .C2(G162gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1347gat));
  NOR2_X1   g616(.A1(new_n590_), .A2(new_n494_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n540_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n779_), .A2(new_n361_), .A3(new_n568_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G169gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n392_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n824_), .B(new_n825_), .C1(new_n826_), .C2(new_n821_), .ZN(G1348gat));
  AOI21_X1  g626(.A(new_n362_), .B1(new_n741_), .B2(new_n772_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(G176gat), .A3(new_n313_), .A4(new_n820_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n830_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n779_), .A2(new_n820_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n313_), .A3(new_n361_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n831_), .A2(new_n832_), .B1(new_n834_), .B2(new_n393_), .ZN(G1349gat));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n361_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n583_), .A2(new_n430_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n828_), .A2(new_n285_), .A3(new_n820_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n836_), .A2(new_n837_), .B1(new_n396_), .B2(new_n838_), .ZN(G1350gat));
  NAND4_X1  g638(.A1(new_n779_), .A2(new_n616_), .A3(new_n361_), .A4(new_n820_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G190gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n582_), .B1(new_n437_), .B2(new_n434_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT125), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n779_), .A2(new_n361_), .A3(new_n820_), .A4(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT126), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n841_), .A2(new_n847_), .A3(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1351gat));
  NOR2_X1   g648(.A1(new_n819_), .A2(new_n361_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n801_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n569_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n342_), .ZN(G1352gat));
  INV_X1    g652(.A(new_n851_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n313_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g655(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n801_), .A2(new_n285_), .A3(new_n850_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n859_), .A2(KEYINPUT127), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT127), .B1(new_n859_), .B2(new_n861_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n857_), .B1(new_n851_), .B2(new_n583_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(G1354gat));
  AND3_X1   g664(.A1(new_n854_), .A2(G218gat), .A3(new_n616_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G218gat), .B1(new_n854_), .B2(new_n582_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1355gat));
endmodule


