//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT10), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n221_), .B2(KEYINPUT9), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n211_), .A2(new_n213_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT65), .B1(new_n219_), .B2(new_n220_), .ZN(new_n225_));
  INV_X1    g024(.A(G85gat), .ZN(new_n226_));
  INV_X1    g025(.A(G92gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n212_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n204_), .A3(new_n203_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n216_), .A3(new_n217_), .A4(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n224_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n231_), .A2(new_n224_), .A3(new_n235_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n223_), .B(KEYINPUT69), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT65), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n229_), .B1(new_n228_), .B2(new_n212_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n235_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n231_), .A2(new_n224_), .A3(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT69), .B1(new_n245_), .B2(new_n223_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G43gat), .B(G50gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT15), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n223_), .B(KEYINPUT66), .C1(new_n236_), .C2(new_n237_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT66), .B1(new_n245_), .B2(new_n223_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n250_), .B(new_n251_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT35), .Z(new_n262_));
  NAND4_X1  g061(.A1(new_n254_), .A2(new_n258_), .A3(new_n259_), .A4(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n258_), .B(new_n262_), .C1(new_n247_), .C2(new_n253_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT75), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT35), .A3(new_n261_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G190gat), .B(G218gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(G134gat), .B(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT36), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT74), .Z(new_n276_));
  NAND4_X1  g075(.A1(new_n265_), .A2(new_n263_), .A3(new_n267_), .A4(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(KEYINPUT76), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(KEYINPUT76), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n202_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT77), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n268_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n265_), .A2(new_n263_), .A3(new_n267_), .A4(KEYINPUT77), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n272_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT37), .B1(new_n285_), .B2(new_n277_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT78), .B1(new_n280_), .B2(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G127gat), .B(G155gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G211gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT16), .B(G183gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G57gat), .B(G64gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G78gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(G78gat), .B1(new_n305_), .B2(new_n300_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n306_), .A3(KEYINPUT11), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n299_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n299_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT80), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n314_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G1gat), .A2(G8gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT14), .ZN(new_n319_));
  INV_X1    g118(.A(G15gat), .ZN(new_n320_));
  INV_X1    g119(.A(G22gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G15gat), .A2(G22gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n324_), .A2(KEYINPUT79), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(KEYINPUT79), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G1gat), .B(G8gat), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n317_), .B(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(KEYINPUT17), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n297_), .B1(new_n332_), .B2(new_n295_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n331_), .A2(KEYINPUT81), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n291_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339_));
  NOR3_X1   g138(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  AOI211_X1 g145(.A(new_n340_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n348_), .B(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n352_), .B2(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n349_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n352_), .B2(new_n349_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT22), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT22), .B1(new_n358_), .B2(new_n359_), .ZN(new_n361_));
  INV_X1    g160(.A(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n356_), .A2(new_n357_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n354_), .B1(new_n342_), .B2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G211gat), .B(G218gat), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G197gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n368_), .A2(G204gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(G204gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT21), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n368_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n370_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n367_), .B(new_n371_), .C1(new_n374_), .C2(KEYINPUT21), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT21), .A3(new_n366_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n365_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n353_), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G169gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n342_), .B1(new_n385_), .B2(new_n362_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n356_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n347_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n377_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT95), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n393_), .A3(new_n377_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n380_), .A2(new_n383_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n365_), .A2(new_n377_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(KEYINPUT20), .C1(new_n390_), .C2(new_n377_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n383_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT18), .B(G64gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n380_), .A2(new_n398_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(new_n383_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n404_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n410_), .A3(KEYINPUT99), .ZN(new_n411_));
  AOI211_X1 g210(.A(KEYINPUT99), .B(new_n404_), .C1(new_n395_), .C2(new_n399_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n339_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n409_), .A2(new_n404_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n339_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  INV_X1    g220(.A(G134gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT89), .B(G127gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G155gat), .B(G162gat), .Z(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT90), .A2(KEYINPUT2), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT90), .A2(KEYINPUT2), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n432_), .B(new_n433_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n428_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT1), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n428_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n427_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n436_), .B(new_n441_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT4), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n427_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n420_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n444_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n449_), .A2(new_n420_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n226_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT0), .B(G57gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n452_), .B(new_n453_), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OR3_X1    g254(.A1(new_n448_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n427_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT88), .B(KEYINPUT30), .Z(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G15gat), .B(G43gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT31), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G99gat), .Z(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n365_), .B(new_n467_), .ZN(new_n468_));
  OR3_X1    g267(.A1(new_n462_), .A2(new_n463_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT28), .B(G22gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n442_), .A2(KEYINPUT29), .ZN(new_n474_));
  INV_X1    g273(.A(G50gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n474_), .A2(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n473_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n481_), .A3(KEYINPUT93), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n442_), .A2(KEYINPUT29), .B1(new_n375_), .B2(new_n376_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G78gat), .B(G106gat), .Z(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n481_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT91), .B1(new_n485_), .B2(new_n486_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n488_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n486_), .B1(new_n485_), .B2(KEYINPUT93), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n493_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n471_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n419_), .A2(KEYINPUT100), .A3(new_n458_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT100), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT99), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n416_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n412_), .B1(new_n501_), .B2(new_n406_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n458_), .B(new_n417_), .C1(new_n502_), .C2(new_n339_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n503_), .B2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n456_), .A2(new_n457_), .B1(new_n409_), .B2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT97), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT97), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT98), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n492_), .A2(new_n495_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n454_), .B1(new_n449_), .B2(new_n420_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n445_), .A2(new_n420_), .A3(new_n447_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT96), .B(new_n454_), .C1(new_n449_), .C2(new_n420_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n415_), .A2(new_n521_), .A3(new_n416_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n457_), .B(KEYINPUT33), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n507_), .A2(new_n509_), .A3(KEYINPUT98), .A4(new_n510_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n513_), .A2(new_n515_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n503_), .A2(new_n514_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n471_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n505_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n309_), .A2(new_n310_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n298_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n312_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n223_), .B1(new_n237_), .B2(new_n236_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n538_), .B2(new_n255_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT68), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n255_), .A3(new_n535_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n532_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT12), .B1(new_n311_), .B2(new_n313_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n247_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n536_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n238_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n545_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT70), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n546_), .A2(new_n551_), .B1(new_n541_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n539_), .B2(new_n532_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n314_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(KEYINPUT72), .A3(new_n531_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n543_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT5), .B(G176gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n543_), .A2(new_n559_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n569_), .B2(KEYINPUT13), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n330_), .A2(new_n253_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT84), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n252_), .B(KEYINPUT82), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n330_), .A2(KEYINPUT83), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT83), .B1(new_n330_), .B2(new_n578_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n575_), .B(new_n577_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n330_), .A2(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n330_), .A2(new_n578_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT83), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n583_), .B1(new_n586_), .B2(new_n579_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n587_), .B2(new_n576_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G169gat), .B(G197gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT85), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n588_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n574_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n530_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n338_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n458_), .B(KEYINPUT101), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n601_), .A2(new_n602_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(KEYINPUT103), .A3(new_n602_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n285_), .A2(new_n277_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n596_), .A2(new_n335_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(KEYINPUT102), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(KEYINPUT102), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n608_), .B(new_n530_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n458_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .A4(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT104), .Z(G1324gat));
  NAND2_X1  g414(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n616_));
  OAI211_X1 g415(.A(G8gat), .B(new_n616_), .C1(new_n612_), .C2(new_n419_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G8gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n419_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n598_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n619_), .A2(new_n622_), .A3(new_n623_), .A4(new_n625_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n612_), .B2(new_n528_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT41), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n598_), .A2(new_n320_), .A3(new_n471_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n612_), .B2(new_n515_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n598_), .A2(new_n321_), .A3(new_n514_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  NOR3_X1   g436(.A1(new_n574_), .A2(new_n335_), .A3(new_n595_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n530_), .A2(new_n639_), .A3(new_n291_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n530_), .B2(new_n291_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI221_X1 g443(.A(new_n638_), .B1(KEYINPUT107), .B2(KEYINPUT44), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G29gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n600_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n335_), .A2(new_n608_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n530_), .A2(new_n596_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n458_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n649_), .A2(new_n654_), .ZN(G1328gat));
  OAI21_X1  g454(.A(G36gat), .B1(new_n646_), .B2(new_n419_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n621_), .A2(KEYINPUT108), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n621_), .A2(KEYINPUT108), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n651_), .A2(G36gat), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n656_), .A2(new_n658_), .A3(new_n664_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n657_), .A2(KEYINPUT109), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1329gat));
  AOI21_X1  g466(.A(G43gat), .B1(new_n652_), .B2(new_n471_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n471_), .A2(G43gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n644_), .A2(new_n645_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n644_), .A2(new_n645_), .A3(KEYINPUT110), .A4(new_n669_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n674_), .B(new_n676_), .ZN(G1330gat));
  OAI21_X1  g476(.A(G50gat), .B1(new_n646_), .B2(new_n515_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n514_), .A2(new_n475_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT112), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n651_), .B2(new_n680_), .ZN(G1331gat));
  AOI21_X1  g480(.A(new_n594_), .B1(new_n505_), .B2(new_n529_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT113), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT113), .B(new_n594_), .C1(new_n505_), .C2(new_n529_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n684_), .A2(new_n338_), .A3(new_n685_), .A4(new_n573_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n600_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n682_), .A2(new_n608_), .A3(new_n335_), .A4(new_n574_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT114), .Z(new_n689_));
  AND2_X1   g488(.A1(new_n653_), .A2(G57gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n661_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n686_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n686_), .A2(new_n700_), .A3(new_n471_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n689_), .A2(new_n471_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G71gat), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1334gat));
  NAND3_X1  g505(.A1(new_n686_), .A2(new_n302_), .A3(new_n514_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n689_), .A2(new_n514_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G78gat), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1335gat));
  OR2_X1    g511(.A1(new_n682_), .A2(new_n683_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n682_), .A2(new_n683_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n574_), .A3(new_n650_), .A4(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT116), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n684_), .A2(new_n685_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT116), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n574_), .A4(new_n650_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n600_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n574_), .A2(new_n336_), .A3(new_n595_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT117), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT118), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n723_), .B(KEYINPUT118), .C1(new_n641_), .C2(new_n640_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n458_), .A2(new_n226_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n721_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n720_), .B2(new_n621_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n661_), .A2(new_n227_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n728_), .B2(new_n732_), .ZN(G1337gat));
  NOR2_X1   g532(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n734_));
  AND2_X1   g533(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n209_), .A2(new_n210_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n736_), .A3(new_n471_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n726_), .A2(new_n471_), .A3(new_n727_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G99gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n734_), .B(new_n735_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n740_));
  AND4_X1   g539(.A1(KEYINPUT119), .A2(new_n737_), .A3(KEYINPUT51), .A4(new_n739_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n720_), .A2(new_n203_), .A3(new_n514_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n724_), .A2(new_n515_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G106gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G106gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n743_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  NOR3_X1   g551(.A1(new_n648_), .A2(new_n621_), .A3(new_n496_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n337_), .A2(new_n595_), .A3(new_n573_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT54), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n337_), .A2(new_n757_), .A3(new_n595_), .A4(new_n573_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n582_), .B(new_n591_), .C1(new_n587_), .C2(new_n576_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n575_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n577_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI221_X1 g564(.A(new_n577_), .B1(new_n330_), .B2(new_n578_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n591_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n762_), .A2(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n568_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n539_), .A2(new_n554_), .A3(new_n532_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT72), .B1(new_n556_), .B2(new_n531_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n541_), .A2(new_n552_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n544_), .B(new_n545_), .C1(new_n548_), .C2(new_n238_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT70), .B1(new_n549_), .B2(new_n550_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n770_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n532_), .B1(new_n777_), .B2(new_n540_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n558_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n564_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n781_), .C2(new_n564_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n594_), .A2(new_n567_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n769_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n608_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n760_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n768_), .A2(new_n567_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT121), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n768_), .A2(new_n795_), .A3(new_n567_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n564_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n782_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT122), .B(KEYINPUT56), .C1(new_n781_), .C2(new_n564_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n797_), .B(KEYINPUT58), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n291_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n792_), .A2(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n790_), .A2(new_n760_), .A3(new_n791_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n336_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n754_), .B1(new_n759_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n594_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n808_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n792_), .A2(new_n806_), .A3(KEYINPUT123), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n335_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n759_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n753_), .A2(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n817_), .A2(new_n819_), .B1(new_n818_), .B2(new_n810_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n594_), .A2(G113gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n811_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n820_), .B2(new_n573_), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n825_), .A2(KEYINPUT60), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT124), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(G1341gat));
  AOI21_X1  g629(.A(G127gat), .B1(new_n810_), .B2(new_n335_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n335_), .A2(G127gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n821_), .B2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n810_), .B2(new_n791_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n291_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n422_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n821_), .B2(new_n836_), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n759_), .A2(new_n809_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n515_), .A2(new_n471_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n693_), .A2(new_n648_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n594_), .A3(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT125), .B(G141gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1344gat));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n574_), .A3(new_n842_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT126), .B(G148gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n335_), .A3(new_n842_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  NOR3_X1   g650(.A1(new_n840_), .A2(new_n648_), .A3(new_n693_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n791_), .ZN(new_n853_));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n835_), .A2(new_n854_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n853_), .A2(new_n854_), .B1(new_n852_), .B2(new_n855_), .ZN(G1347gat));
  NOR3_X1   g655(.A1(new_n661_), .A2(new_n600_), .A3(new_n496_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n594_), .B(new_n857_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G169gat), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n792_), .A2(new_n806_), .A3(KEYINPUT123), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT123), .B1(new_n792_), .B2(new_n806_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n808_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n759_), .B1(new_n862_), .B2(new_n335_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n594_), .A3(new_n385_), .A4(new_n857_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1348gat));
  NAND4_X1  g668(.A1(new_n863_), .A2(new_n362_), .A3(new_n574_), .A4(new_n857_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n838_), .A2(new_n574_), .A3(new_n857_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n362_), .ZN(G1349gat));
  NAND3_X1  g671(.A1(new_n816_), .A2(new_n335_), .A3(new_n857_), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n345_), .B(G183gat), .S(new_n873_), .Z(G1350gat));
  OAI211_X1 g673(.A(new_n291_), .B(new_n857_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G190gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n863_), .A2(new_n791_), .A3(new_n346_), .A4(new_n857_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n877_), .A3(KEYINPUT127), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  NOR3_X1   g681(.A1(new_n840_), .A2(new_n653_), .A3(new_n661_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n594_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G197gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n368_), .A3(new_n594_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1352gat));
  NOR2_X1   g686(.A1(new_n661_), .A2(new_n653_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n841_), .A2(new_n574_), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  AND2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n883_), .B(new_n335_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n883_), .A2(new_n335_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n891_), .ZN(G1354gat));
  NAND2_X1  g694(.A1(new_n883_), .A2(new_n791_), .ZN(new_n896_));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n835_), .A2(new_n897_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n896_), .A2(new_n897_), .B1(new_n883_), .B2(new_n898_), .ZN(G1355gat));
endmodule


