//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_;
  XOR2_X1   g000(.A(G176gat), .B(G204gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G230gat), .A2(G233gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n210_), .A2(new_n211_), .B1(new_n213_), .B2(KEYINPUT66), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n209_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n214_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(KEYINPUT67), .C1(new_n221_), .C2(new_n212_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G85gat), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G92gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n210_), .A2(KEYINPUT10), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n210_), .A2(KEYINPUT10), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(KEYINPUT64), .A3(new_n211_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n211_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n225_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G92gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n230_), .A2(new_n232_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT9), .B1(new_n230_), .B2(new_n232_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT65), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n231_), .A2(G92gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n229_), .A2(G85gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n230_), .A2(new_n232_), .A3(new_n243_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n238_), .B(new_n241_), .C1(new_n246_), .C2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n220_), .B1(new_n221_), .B2(new_n212_), .ZN(new_n254_));
  OAI22_X1  g053(.A1(new_n254_), .A2(new_n225_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n228_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n234_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G57gat), .B(G64gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n260_));
  XOR2_X1   g059(.A(G71gat), .B(G78gat), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n257_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n234_), .A2(new_n253_), .A3(new_n256_), .A4(new_n264_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(new_n269_), .A3(new_n265_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n208_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n207_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n206_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n206_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n274_), .A2(KEYINPUT69), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n274_), .B2(new_n275_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT70), .B(G43gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  INV_X1    g083(.A(G50gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n283_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT74), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n298_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n291_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n293_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(new_n290_), .A3(new_n289_), .A4(new_n300_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n282_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n300_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n289_), .A2(KEYINPUT15), .A3(new_n290_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT15), .B1(new_n289_), .B2(new_n290_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n282_), .A3(new_n306_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n281_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n324_));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G64gat), .B(G92gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  INV_X1    g132(.A(G183gat), .ZN(new_n334_));
  INV_X1    g133(.A(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT23), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT88), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(KEYINPUT88), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n341_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n350_), .B2(new_n349_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT25), .B(G183gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n335_), .A2(KEYINPUT26), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n335_), .A2(KEYINPUT26), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n338_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n336_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n348_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G197gat), .B(G204gat), .Z(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n333_), .B1(new_n362_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(G183gat), .B2(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n360_), .B(KEYINPUT80), .C1(G183gat), .C2(G190gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n344_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n354_), .B1(new_n355_), .B2(KEYINPUT78), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n355_), .A2(KEYINPUT78), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n353_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n352_), .B(new_n339_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n369_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n332_), .B1(new_n370_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT20), .B(new_n332_), .C1(new_n362_), .C2(new_n369_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n329_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n381_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n346_), .A2(new_n347_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n380_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n331_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI211_X1 g189(.A(new_n333_), .B(new_n331_), .C1(new_n388_), .C2(new_n380_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n384_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n393_), .A3(new_n328_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n386_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT94), .A4(new_n328_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n370_), .A2(new_n332_), .A3(new_n381_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n380_), .A2(new_n361_), .A3(new_n345_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT20), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n331_), .B1(new_n384_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n329_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n396_), .B1(new_n406_), .B2(KEYINPUT27), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(new_n231_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT0), .B(G57gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G141gat), .A2(G148gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT82), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT2), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419_));
  OR4_X1    g218(.A1(new_n419_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n416_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n421_), .A2(KEYINPUT2), .B1(new_n419_), .B2(KEYINPUT3), .ZN(new_n422_));
  INV_X1    g221(.A(G141gat), .ZN(new_n423_));
  INV_X1    g222(.A(G148gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n419_), .B2(KEYINPUT3), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n420_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n414_), .B(new_n415_), .C1(new_n418_), .C2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G127gat), .B(G134gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G120gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n417_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n414_), .A2(KEYINPUT1), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n414_), .A2(KEYINPUT1), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n415_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n425_), .A2(KEYINPUT83), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n425_), .A2(KEYINPUT83), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n428_), .A2(new_n431_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n431_), .B(KEYINPUT81), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n428_), .A2(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n413_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(KEYINPUT4), .A3(new_n443_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n441_), .A2(new_n442_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT90), .B(KEYINPUT4), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n411_), .B(new_n445_), .C1(new_n450_), .C2(new_n412_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n411_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n412_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n453_), .B2(new_n444_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G78gat), .B(G106gat), .Z(new_n456_));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n428_), .A2(new_n438_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n369_), .B(new_n457_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(KEYINPUT29), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n428_), .B2(new_n438_), .ZN(new_n462_));
  OAI211_X1 g261(.A(G228gat), .B(G233gat), .C1(new_n462_), .C2(new_n380_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(KEYINPUT87), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n463_), .A3(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  INV_X1    g267(.A(new_n466_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n464_), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n442_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT28), .B1(new_n442_), .B2(KEYINPUT29), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G22gat), .B(G50gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n469_), .B1(KEYINPUT87), .B2(new_n464_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n467_), .A2(new_n470_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT85), .B1(new_n469_), .B2(new_n464_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n455_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT95), .B1(new_n407_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n455_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n394_), .A2(new_n397_), .B1(new_n404_), .B2(new_n329_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n395_), .B1(new_n485_), .B2(new_n399_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n483_), .B(new_n484_), .C1(new_n486_), .C2(new_n396_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n451_), .A2(new_n454_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n328_), .A2(KEYINPUT32), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n390_), .A2(new_n393_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT93), .A4(new_n489_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n404_), .A2(KEYINPUT32), .A3(new_n328_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n488_), .A2(new_n492_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n454_), .B(new_n496_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n447_), .A2(KEYINPUT91), .A3(new_n439_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT91), .B1(new_n447_), .B2(new_n439_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n413_), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n446_), .A2(new_n449_), .A3(new_n412_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT92), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n502_), .A3(new_n411_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(KEYINPUT92), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n394_), .B(new_n386_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n495_), .B1(new_n497_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n478_), .A2(new_n480_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n482_), .A2(new_n487_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n375_), .A2(new_n379_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G227gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(new_n441_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT30), .B(G15gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G43gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n513_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n509_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n507_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT96), .B1(new_n407_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n524_), .B(new_n507_), .C1(new_n486_), .C2(new_n396_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n523_), .A2(new_n525_), .A3(new_n455_), .A4(new_n519_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n323_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n309_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n264_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT77), .Z(new_n539_));
  NOR2_X1   g338(.A1(new_n530_), .A2(new_n536_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT76), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n257_), .A2(new_n291_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n257_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(KEYINPUT35), .A3(new_n546_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G134gat), .B(G162gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n543_), .A2(new_n544_), .A3(new_n557_), .A4(new_n547_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT73), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n549_), .A2(new_n561_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n564_));
  INV_X1    g363(.A(new_n549_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n558_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(KEYINPUT37), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n542_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n527_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n295_), .A3(new_n488_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n568_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n542_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n527_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n578_), .B2(new_n455_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n574_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n579_), .A3(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(new_n407_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(G8gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n527_), .A2(new_n407_), .A3(new_n577_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(G8gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n587_), .B2(G8gat), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(G1325gat));
  OAI21_X1  g394(.A(G15gat), .B1(new_n578_), .B2(new_n520_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT41), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT41), .ZN(new_n598_));
  INV_X1    g397(.A(G15gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n572_), .A2(new_n599_), .A3(new_n519_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n507_), .B(KEYINPUT99), .Z(new_n603_));
  NAND3_X1  g402(.A1(new_n572_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G22gat), .B1(new_n578_), .B2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT42), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT42), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT100), .ZN(G1327gat));
  NAND3_X1  g409(.A1(new_n281_), .A2(new_n322_), .A3(new_n542_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT101), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n521_), .A2(new_n526_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n569_), .A2(new_n570_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n569_), .A2(new_n570_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT43), .B(new_n617_), .C1(new_n521_), .C2(new_n526_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n612_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT44), .B(new_n612_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n488_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G29gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n542_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n568_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n527_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n455_), .A2(G29gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT46), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n621_), .A2(new_n407_), .A3(new_n622_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G36gat), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n582_), .A2(G36gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n527_), .A2(new_n626_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n527_), .A2(new_n626_), .A3(new_n636_), .A4(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n630_), .A2(new_n631_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n633_), .B1(new_n635_), .B2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n632_), .B(new_n645_), .C1(new_n634_), .C2(G36gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1329gat));
  NAND4_X1  g448(.A1(new_n621_), .A2(G43gat), .A3(new_n519_), .A4(new_n622_), .ZN(new_n650_));
  INV_X1    g449(.A(G43gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n627_), .B2(new_n520_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1330gat));
  NAND3_X1  g454(.A1(new_n621_), .A2(new_n522_), .A3(new_n622_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n285_), .B1(new_n656_), .B2(KEYINPUT106), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(KEYINPUT106), .B2(new_n656_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n527_), .A2(new_n285_), .A3(new_n603_), .A4(new_n626_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1331gat));
  AOI211_X1 g459(.A(new_n322_), .B(new_n281_), .C1(new_n521_), .C2(new_n526_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n577_), .ZN(new_n662_));
  INV_X1    g461(.A(G57gat), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n455_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT109), .ZN(new_n665_));
  INV_X1    g464(.A(new_n281_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT107), .B1(new_n571_), .B2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n322_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n571_), .A2(new_n666_), .A3(KEYINPUT107), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n614_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT108), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT108), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n488_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n665_), .B1(new_n663_), .B2(new_n674_), .ZN(G1332gat));
  OAI21_X1  g474(.A(G64gat), .B1(new_n662_), .B2(new_n582_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT48), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n582_), .A2(G64gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n670_), .B2(new_n678_), .ZN(G1333gat));
  OR3_X1    g478(.A1(new_n670_), .A2(G71gat), .A3(new_n520_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n661_), .A2(new_n519_), .A3(new_n577_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G71gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT110), .Z(G1334gat));
  OR3_X1    g485(.A1(new_n670_), .A2(G78gat), .A3(new_n605_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G78gat), .B1(new_n662_), .B2(new_n605_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT50), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT50), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT111), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(new_n687_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1335gat));
  AND2_X1   g494(.A1(new_n661_), .A2(new_n626_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n488_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT112), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n616_), .A2(new_n618_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n281_), .A2(new_n625_), .A3(new_n322_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n231_), .A3(new_n455_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1336gat));
  AOI21_X1  g502(.A(G92gat), .B1(new_n696_), .B2(new_n407_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n582_), .A2(new_n229_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1337gat));
  OAI21_X1  g506(.A(G99gat), .B1(new_n701_), .B2(new_n520_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n661_), .A2(new_n237_), .A3(new_n519_), .A4(new_n626_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT113), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT51), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n711_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n708_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n696_), .A2(new_n211_), .A3(new_n522_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n522_), .B(new_n700_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G106gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G106gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g522(.A1(new_n523_), .A2(new_n525_), .A3(new_n488_), .A4(new_n519_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT120), .Z(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT58), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n268_), .A2(new_n208_), .A3(new_n270_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT55), .ZN(new_n729_));
  INV_X1    g528(.A(new_n271_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n268_), .A2(new_n270_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(KEYINPUT55), .A3(new_n207_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n271_), .A2(KEYINPUT114), .A3(KEYINPUT55), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n206_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(KEYINPUT117), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n206_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT117), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n277_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n274_), .A2(KEYINPUT69), .A3(new_n275_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n306_), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n305_), .A2(new_n300_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n282_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n316_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n282_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT115), .B1(new_n752_), .B2(new_n317_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n312_), .A2(new_n751_), .A3(new_n306_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n318_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n318_), .A3(KEYINPUT116), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n744_), .A2(new_n745_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n743_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n727_), .B1(new_n740_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n741_), .A2(new_n742_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(KEYINPUT58), .A3(new_n743_), .A4(new_n760_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n615_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n762_), .A2(new_n615_), .A3(new_n767_), .A4(KEYINPUT118), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n322_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n758_), .A2(new_n759_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n278_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n568_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n568_), .C1(new_n774_), .C2(new_n777_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT119), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n321_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n576_), .B1(new_n785_), .B2(new_n776_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n780_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n542_), .B1(new_n772_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n322_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n571_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n571_), .B2(new_n790_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n726_), .B1(new_n789_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G113gat), .B1(new_n796_), .B2(new_n322_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n768_), .A2(new_n780_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n781_), .A2(KEYINPUT119), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n783_), .A3(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n625_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n798_), .B(new_n725_), .C1(new_n803_), .C2(new_n794_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT121), .B(new_n804_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n322_), .A2(G113gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT122), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n797_), .B1(new_n809_), .B2(new_n811_), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n796_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n813_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n666_), .B(new_n804_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n816_), .A2(KEYINPUT123), .ZN(new_n817_));
  OAI21_X1  g616(.A(G120gat), .B1(new_n816_), .B2(KEYINPUT123), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n817_), .B2(new_n818_), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n796_), .B2(new_n625_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n625_), .A2(G127gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n809_), .B2(new_n821_), .ZN(G1342gat));
  NAND4_X1  g621(.A1(new_n770_), .A2(new_n802_), .A3(new_n780_), .A4(new_n771_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n794_), .B1(new_n823_), .B2(new_n542_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(new_n568_), .A3(new_n726_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT124), .B1(new_n825_), .B2(G134gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n789_), .A2(new_n795_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n576_), .A3(new_n725_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829_));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n617_), .A2(new_n830_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n809_), .B2(new_n833_), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n520_), .A2(new_n522_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n824_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n407_), .A2(new_n455_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n423_), .A3(new_n322_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G141gat), .B1(new_n838_), .B2(new_n321_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1344gat));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n424_), .A3(new_n666_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G148gat), .B1(new_n838_), .B2(new_n281_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1345gat));
  NAND3_X1  g644(.A1(new_n836_), .A2(new_n625_), .A3(new_n837_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n838_), .A2(new_n849_), .A3(new_n617_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n839_), .A2(new_n576_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n849_), .B2(new_n851_), .ZN(G1347gat));
  OR2_X1    g651(.A1(new_n803_), .A2(new_n794_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n582_), .A2(new_n488_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n519_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n603_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G169gat), .B1(new_n857_), .B2(new_n321_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT62), .B(G169gat), .C1(new_n857_), .C2(new_n321_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n857_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n322_), .A3(new_n342_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n861_), .A3(new_n863_), .ZN(G1348gat));
  AOI21_X1  g663(.A(G176gat), .B1(new_n862_), .B2(new_n666_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n824_), .A2(new_n522_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n855_), .A2(new_n343_), .A3(new_n281_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1349gat));
  INV_X1    g667(.A(new_n353_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n853_), .A2(new_n869_), .A3(new_n625_), .A4(new_n856_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n855_), .A2(new_n542_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n866_), .A2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT125), .B(new_n870_), .C1(new_n872_), .C2(G183gat), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  INV_X1    g673(.A(new_n870_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G183gat), .B1(new_n866_), .B2(new_n871_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(G1350gat));
  NAND4_X1  g677(.A1(new_n862_), .A2(new_n354_), .A3(new_n355_), .A4(new_n576_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n862_), .A2(new_n615_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n881_), .B2(new_n335_), .ZN(G1351gat));
  NAND3_X1  g681(.A1(new_n836_), .A2(new_n322_), .A3(new_n854_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g683(.A1(new_n836_), .A2(new_n666_), .A3(new_n854_), .ZN(new_n885_));
  INV_X1    g684(.A(G204gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1353gat));
  AND2_X1   g686(.A1(new_n836_), .A2(new_n854_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n542_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n888_), .A2(new_n892_), .A3(new_n889_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1354gat));
  NAND2_X1  g695(.A1(new_n888_), .A2(new_n576_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT127), .B(G218gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n617_), .A2(new_n899_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n897_), .A2(new_n899_), .B1(new_n888_), .B2(new_n900_), .ZN(G1355gat));
endmodule


