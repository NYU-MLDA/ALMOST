//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT85), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT30), .B(G15gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT31), .Z(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT23), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT81), .B1(new_n224_), .B2(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n223_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT81), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n222_), .A3(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n218_), .A2(new_n219_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT83), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n221_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n214_), .B(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n236_), .A2(new_n213_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n237_));
  OAI22_X1  g036(.A1(new_n228_), .A2(new_n229_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n210_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n210_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n249_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n251_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n255_), .A3(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT88), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT3), .ZN(new_n265_));
  OR3_X1    g064(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n266_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n262_), .B(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n264_), .B(new_n267_), .C1(new_n274_), .C2(new_n261_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT29), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n247_), .B(new_n248_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n278_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT89), .B1(new_n281_), .B2(KEYINPUT87), .ZN(new_n282_));
  OAI211_X1 g081(.A(G228gat), .B(G233gat), .C1(new_n278_), .C2(new_n247_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G78gat), .B(G106gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n272_), .A2(new_n289_), .A3(new_n275_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT28), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n290_), .A2(KEYINPUT28), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n288_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n291_), .A3(new_n287_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT90), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n285_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n280_), .B(new_n302_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n286_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n300_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n286_), .B2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n205_), .A2(new_n276_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT93), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n202_), .B(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(new_n204_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n204_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n275_), .B(new_n272_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n309_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n205_), .A2(KEYINPUT93), .A3(new_n276_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT4), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT94), .Z(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT95), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n309_), .A2(KEYINPUT4), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n321_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  INV_X1    g128(.A(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n328_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT33), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n326_), .A2(new_n337_), .A3(new_n328_), .A4(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n236_), .A2(new_n213_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n226_), .A2(new_n223_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n340_), .A2(new_n217_), .A3(new_n222_), .A4(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n221_), .A3(new_n232_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(new_n258_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n238_), .A2(new_n258_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND4_X1   g149(.A1(KEYINPUT20), .A2(new_n346_), .A3(new_n347_), .A4(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n258_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT91), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n345_), .A2(KEYINPUT92), .A3(new_n258_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT92), .B1(new_n345_), .B2(new_n258_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n357_), .B(KEYINPUT20), .C1(new_n238_), .C2(new_n258_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n359_), .B2(new_n349_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  INV_X1    g160(.A(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT18), .B(G64gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n319_), .A2(new_n327_), .A3(new_n325_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n334_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n366_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n339_), .A2(new_n368_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n375_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n328_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n333_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n335_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT96), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n349_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n359_), .B2(new_n349_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n380_), .A3(new_n349_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n360_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n379_), .B(new_n386_), .C1(new_n384_), .C2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n308_), .B1(new_n373_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n286_), .A2(new_n303_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n300_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n286_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n379_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n365_), .B(new_n351_), .C1(new_n359_), .C2(new_n349_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n367_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n383_), .A2(new_n365_), .A3(new_n385_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT27), .A3(new_n372_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n393_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n246_), .B1(new_n389_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n307_), .A3(new_n399_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n379_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n397_), .A2(new_n307_), .A3(new_n399_), .A4(KEYINPUT98), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n245_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n401_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT67), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT66), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT66), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT6), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n414_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n412_), .A2(KEYINPUT6), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n410_), .A2(KEYINPUT66), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT67), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n417_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G85gat), .B(G92gat), .Z(new_n429_));
  INV_X1    g228(.A(KEYINPUT8), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n429_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT8), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT10), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT64), .B(G106gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT65), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n330_), .A2(new_n362_), .A3(KEYINPUT9), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n429_), .B2(KEYINPUT9), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n417_), .A2(new_n423_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n436_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G64gat), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n451_));
  XOR2_X1   g250(.A(G71gat), .B(G78gat), .Z(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n448_), .A2(KEYINPUT68), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G230gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n428_), .A2(new_n431_), .B1(new_n434_), .B2(KEYINPUT8), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n445_), .A2(new_n446_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n436_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT68), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT12), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n448_), .A2(new_n467_), .A3(new_n456_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT69), .B1(new_n469_), .B2(new_n458_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT69), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n471_), .B(new_n459_), .C1(new_n466_), .C2(new_n468_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n465_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G120gat), .B(G148gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G204gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT5), .B(G176gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n465_), .B(new_n477_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n479_), .A2(KEYINPUT13), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT13), .B1(new_n479_), .B2(new_n480_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT75), .B(G15gat), .ZN(new_n486_));
  INV_X1    g285(.A(G22gat), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT76), .B(G1gat), .ZN(new_n489_));
  INV_X1    g288(.A(G8gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n487_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G43gat), .B(G50gat), .Z(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT15), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n505_), .B(KEYINPUT80), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n498_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n498_), .B(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G169gat), .B(G197gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n515_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n485_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n408_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n506_), .B1(new_n436_), .B2(new_n447_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n505_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n460_), .A2(new_n461_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n505_), .B(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n533_), .B2(KEYINPUT70), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n526_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT35), .B(new_n528_), .C1(new_n523_), .C2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n533_), .B1(new_n448_), .B2(new_n505_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G190gat), .B(G218gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT36), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT37), .B1(new_n545_), .B2(KEYINPUT73), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT71), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n529_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n538_), .B1(new_n537_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n526_), .A2(new_n534_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT72), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n535_), .A2(new_n539_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n550_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n545_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n556_), .B2(new_n550_), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT72), .B(new_n549_), .C1(new_n535_), .C2(new_n539_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n560_), .B(new_n544_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n546_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n544_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT74), .ZN(new_n568_));
  INV_X1    g367(.A(new_n546_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n498_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n456_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT78), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT77), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n577_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT17), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT79), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n580_), .A2(KEYINPUT17), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n571_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n522_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n379_), .B(KEYINPUT99), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n489_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n559_), .B(KEYINPUT100), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n586_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n522_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n405_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n597_), .A3(new_n598_), .ZN(G1324gat));
  NAND2_X1  g398(.A1(new_n397_), .A2(new_n399_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n588_), .A2(new_n490_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n600_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(G8gat), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT39), .B(new_n490_), .C1(new_n595_), .C2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n596_), .B2(new_n246_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT41), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT41), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n611_), .B(G15gat), .C1(new_n596_), .C2(new_n246_), .ZN(new_n612_));
  INV_X1    g411(.A(G15gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n588_), .A2(new_n613_), .A3(new_n245_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n610_), .A2(KEYINPUT101), .A3(new_n612_), .A4(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1326gat));
  AOI21_X1  g418(.A(new_n487_), .B1(new_n595_), .B2(new_n308_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n588_), .A2(new_n487_), .A3(new_n308_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1327gat));
  AND3_X1   g422(.A1(new_n568_), .A2(new_n569_), .A3(new_n564_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n569_), .B1(new_n568_), .B2(new_n564_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n571_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n408_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT43), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(KEYINPUT43), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n408_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n634_), .A2(new_n521_), .A3(new_n586_), .A4(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n630_), .A2(KEYINPUT43), .B1(new_n408_), .B2(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n521_), .A2(new_n586_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n589_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G29gat), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n586_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n567_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n522_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n405_), .A2(G29gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  XNOR2_X1  g447(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n637_), .A2(new_n640_), .A3(new_n600_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n600_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n522_), .A2(new_n645_), .A3(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n654_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n649_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n649_), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n660_), .B(new_n657_), .C1(new_n650_), .C2(G36gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1329gat));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n637_), .A2(new_n640_), .A3(new_n245_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G43gat), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n646_), .A2(G43gat), .A3(new_n246_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n663_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT47), .B(new_n666_), .C1(new_n664_), .C2(G43gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1330gat));
  OAI21_X1  g469(.A(G50gat), .B1(new_n641_), .B2(new_n307_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n307_), .A2(G50gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n646_), .B2(new_n673_), .ZN(G1331gat));
  AOI21_X1  g473(.A(new_n519_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n485_), .A3(new_n594_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT109), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(G57gat), .A3(new_n379_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n485_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n408_), .A2(new_n520_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n675_), .A2(KEYINPUT107), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n587_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n686_), .B2(new_n642_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n678_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n688_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g489(.A(new_n686_), .ZN(new_n691_));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n600_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT48), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n677_), .A2(new_n600_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G64gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT48), .B(new_n692_), .C1(new_n677_), .C2(new_n600_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1333gat));
  INV_X1    g497(.A(G71gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n691_), .A2(new_n699_), .A3(new_n245_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n677_), .A2(new_n245_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G71gat), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT49), .B(new_n699_), .C1(new_n677_), .C2(new_n245_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n691_), .A2(new_n706_), .A3(new_n308_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n677_), .A2(new_n308_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G78gat), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT50), .B(new_n706_), .C1(new_n677_), .C2(new_n308_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1335gat));
  AND3_X1   g511(.A1(new_n683_), .A2(new_n645_), .A3(new_n684_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n589_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n715_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n485_), .A2(new_n586_), .A3(new_n520_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n634_), .A2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n330_), .A3(new_n405_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n716_), .A2(new_n717_), .A3(new_n721_), .ZN(G1336gat));
  NOR3_X1   g521(.A1(new_n720_), .A2(new_n362_), .A3(new_n652_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G92gat), .B1(new_n713_), .B2(new_n600_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  NOR2_X1   g524(.A1(new_n246_), .A2(new_n437_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n683_), .A2(new_n645_), .A3(new_n684_), .A4(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n634_), .A2(new_n245_), .A3(new_n719_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n730_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT111), .B1(new_n730_), .B2(G99gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT51), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n729_), .B(new_n735_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1338gat));
  NOR2_X1   g536(.A1(new_n307_), .A2(new_n438_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n713_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n634_), .A2(new_n308_), .A3(new_n719_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n739_), .B(new_n745_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1339gat));
  NAND3_X1  g548(.A1(new_n404_), .A2(new_n245_), .A3(new_n406_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n750_), .A2(new_n642_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT120), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(KEYINPUT59), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n511_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n518_), .B1(new_n512_), .B2(new_n510_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n509_), .A2(new_n513_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n469_), .A2(new_n764_), .A3(KEYINPUT55), .A4(new_n458_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n466_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n469_), .A2(KEYINPUT55), .A3(new_n458_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(KEYINPUT115), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(new_n765_), .A3(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n478_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n480_), .B(new_n761_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n478_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n771_), .A3(new_n770_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(KEYINPUT58), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n478_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n478_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT117), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n782_), .B2(new_n772_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(new_n783_), .A3(new_n571_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n760_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n519_), .A2(new_n480_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n776_), .B2(new_n770_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n567_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n479_), .A2(new_n480_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n786_), .B1(new_n793_), .B2(new_n761_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT116), .B(new_n760_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n788_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n567_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n784_), .A2(new_n792_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n586_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n481_), .A2(new_n483_), .A3(new_n519_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n566_), .A2(new_n644_), .A3(new_n803_), .A4(new_n570_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT114), .B1(new_n804_), .B2(KEYINPUT54), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n626_), .A2(new_n807_), .A3(new_n644_), .A4(new_n803_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n755_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n519_), .A2(G113gat), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n567_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n791_), .B(new_n559_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n644_), .B1(new_n816_), .B2(new_n784_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n809_), .A2(new_n808_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n805_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n751_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n802_), .A2(new_n810_), .A3(KEYINPUT118), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n811_), .B(new_n812_), .C1(new_n823_), .C2(KEYINPUT59), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n820_), .A2(new_n519_), .A3(new_n822_), .A4(new_n821_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(G113gat), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n824_), .A2(new_n828_), .A3(new_n829_), .ZN(G1340gat));
  AOI211_X1 g629(.A(new_n680_), .B(new_n811_), .C1(new_n823_), .C2(KEYINPUT59), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n680_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(KEYINPUT60), .B2(new_n832_), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n831_), .A2(new_n832_), .B1(new_n823_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n820_), .A2(new_n822_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n644_), .A3(new_n821_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n811_), .B1(new_n823_), .B2(KEYINPUT59), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n586_), .A2(new_n836_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n836_), .A2(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n593_), .A3(new_n821_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT121), .B(G134gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n626_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n842_), .A2(new_n843_), .B1(new_n839_), .B2(new_n845_), .ZN(G1343gat));
  NAND4_X1  g645(.A1(new_n652_), .A2(new_n308_), .A3(new_n246_), .A4(new_n589_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT122), .Z(new_n848_));
  NAND3_X1  g647(.A1(new_n837_), .A2(new_n519_), .A3(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g649(.A1(new_n837_), .A2(new_n485_), .A3(new_n848_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g651(.A1(new_n837_), .A2(new_n644_), .A3(new_n848_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  NAND4_X1  g654(.A1(new_n820_), .A2(new_n593_), .A3(new_n822_), .A4(new_n848_), .ZN(new_n856_));
  INV_X1    g655(.A(G162gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n627_), .A2(G162gat), .A3(new_n629_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n820_), .A2(new_n822_), .A3(new_n848_), .A4(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT123), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n863_), .A3(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n308_), .A2(new_n246_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n642_), .A2(new_n866_), .A3(new_n600_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT124), .B1(new_n869_), .B2(new_n520_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n519_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(G169gat), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n870_), .A2(KEYINPUT62), .A3(new_n873_), .A4(G169gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n871_), .A2(new_n519_), .A3(new_n230_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n680_), .A2(new_n231_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n820_), .A2(new_n822_), .A3(new_n868_), .A4(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT125), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT125), .ZN(new_n883_));
  AOI21_X1  g682(.A(G176gat), .B1(new_n871_), .B2(new_n485_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n586_), .A2(new_n223_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n871_), .A2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT126), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n837_), .A2(new_n644_), .A3(new_n868_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n211_), .B2(new_n889_), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n869_), .B2(new_n626_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n871_), .A2(new_n226_), .A3(new_n593_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1351gat));
  AND3_X1   g692(.A1(new_n600_), .A2(new_n393_), .A3(new_n246_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n837_), .A2(new_n519_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g695(.A1(new_n837_), .A2(new_n485_), .A3(new_n894_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g697(.A(new_n586_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT127), .Z(new_n900_));
  NAND3_X1  g699(.A1(new_n837_), .A2(new_n894_), .A3(new_n900_), .ZN(new_n901_));
  OR2_X1    g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1354gat));
  AND2_X1   g702(.A1(new_n837_), .A2(new_n894_), .ZN(new_n904_));
  INV_X1    g703(.A(G218gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n626_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n837_), .A2(new_n593_), .A3(new_n894_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n904_), .A2(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1355gat));
endmodule


