//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_;
  OAI21_X1  g000(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n202_), .B(new_n206_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G85gat), .B(G92gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(new_n212_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n206_), .A2(new_n202_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT8), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n211_), .A2(new_n214_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n216_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT64), .B(G92gat), .Z(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(G85gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n230_));
  INV_X1    g029(.A(new_n220_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT10), .B(G99gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n205_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT15), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT71), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT34), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n243_), .A2(KEYINPUT35), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  AND4_X1   g044(.A1(new_n230_), .A2(new_n229_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(KEYINPUT66), .A2(new_n215_), .B1(new_n222_), .B2(KEYINPUT8), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n225_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n238_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n249_), .B(new_n240_), .C1(KEYINPUT35), .C2(new_n243_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n241_), .A2(new_n240_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G134gat), .B(G162gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT36), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(KEYINPUT36), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n253_), .A2(KEYINPUT72), .A3(new_n257_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT72), .B1(new_n253_), .B2(new_n257_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT37), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n265_));
  XOR2_X1   g064(.A(G71gat), .B(G78gat), .Z(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n266_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT74), .Z(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT73), .B(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n271_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G127gat), .B(G155gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G183gat), .B(G211gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT17), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(KEYINPUT17), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n290_), .B(KEYINPUT76), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n284_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n263_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT78), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n281_), .A2(new_n238_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n281_), .A2(new_n238_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n281_), .A2(KEYINPUT79), .A3(new_n238_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n281_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n304_), .A2(new_n305_), .B1(new_n310_), .B2(new_n239_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n311_), .B2(new_n308_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G113gat), .B(G141gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT80), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT5), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n226_), .A2(new_n234_), .A3(new_n270_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT12), .B1(new_n248_), .B2(new_n270_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n331_));
  INV_X1    g130(.A(new_n270_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n235_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n211_), .A2(new_n214_), .A3(new_n224_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n224_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT8), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n335_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n332_), .B1(new_n339_), .B2(new_n246_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n328_), .B1(new_n340_), .B2(new_n327_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n326_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT67), .ZN(new_n343_));
  INV_X1    g142(.A(new_n328_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n248_), .B2(new_n270_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n331_), .B1(new_n235_), .B2(new_n332_), .ZN(new_n346_));
  AOI211_X1 g145(.A(KEYINPUT12), .B(new_n270_), .C1(new_n226_), .C2(new_n234_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n340_), .A2(new_n327_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n326_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n325_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT68), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n348_), .A2(new_n350_), .A3(KEYINPUT68), .A4(new_n325_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n354_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n362_));
  OAI22_X1  g161(.A1(new_n361_), .A2(new_n362_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n352_), .B1(new_n351_), .B2(new_n326_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT67), .B(new_n325_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n330_), .A2(new_n333_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n341_), .B1(new_n366_), .B2(new_n345_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT68), .B1(new_n367_), .B2(new_n325_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n358_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n364_), .A2(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT69), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n354_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n321_), .B1(new_n363_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT23), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT94), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT25), .B(G183gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT92), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT24), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT93), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(KEYINPUT93), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(G169gat), .B2(G176gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n386_), .B(new_n390_), .C1(new_n393_), .C2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n381_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(new_n391_), .ZN(new_n398_));
  XOR2_X1   g197(.A(KEYINPUT22), .B(G169gat), .Z(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(G176gat), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G204gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n403_), .A2(KEYINPUT90), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(KEYINPUT90), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n402_), .A2(G204gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT21), .ZN(new_n408_));
  XOR2_X1   g207(.A(G211gat), .B(G218gat), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n403_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(KEYINPUT21), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(KEYINPUT21), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n408_), .A2(new_n411_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n379_), .B1(new_n401_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G169gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n417_));
  AOI211_X1 g216(.A(new_n416_), .B(new_n417_), .C1(KEYINPUT83), .C2(KEYINPUT22), .ZN(new_n418_));
  INV_X1    g217(.A(G176gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n398_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT82), .B1(new_n381_), .B2(new_n384_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT81), .B1(new_n425_), .B2(G183gat), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n389_), .B(new_n426_), .C1(new_n387_), .C2(KEYINPUT81), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n428_));
  OAI221_X1 g227(.A(new_n427_), .B1(new_n392_), .B2(new_n382_), .C1(new_n385_), .C2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n414_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n415_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n379_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n430_), .B2(new_n414_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n413_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT95), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT95), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n434_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n433_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT18), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  AND2_X1   g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n441_), .A2(new_n445_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G85gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT0), .B(G57gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G127gat), .B(G134gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT85), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G120gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT89), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT2), .ZN(new_n467_));
  OAI22_X1  g266(.A1(new_n465_), .A2(new_n466_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G155gat), .A2(G162gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT87), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n465_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(KEYINPUT1), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n460_), .B(new_n475_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n459_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n457_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(KEYINPUT4), .A3(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n459_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n453_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n453_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n452_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n452_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(KEYINPUT97), .A3(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n483_), .A2(new_n485_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n496_), .B(new_n497_), .C1(new_n487_), .C2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT33), .B(new_n452_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n445_), .A2(KEYINPUT32), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n441_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n487_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n488_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n493_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n486_), .A2(new_n452_), .A3(new_n488_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n435_), .A2(new_n436_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n434_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT98), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n414_), .B1(new_n401_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n511_), .B2(new_n401_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n432_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n434_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n510_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n517_), .B(new_n379_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n502_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  OAI22_X1  g320(.A1(new_n448_), .A2(new_n501_), .B1(new_n508_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(G78gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n205_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G22gat), .B(G50gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n474_), .A2(new_n529_), .A3(new_n478_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT28), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n413_), .B1(new_n479_), .B2(KEYINPUT29), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n528_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G227gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(G15gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT30), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n430_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n429_), .A2(new_n424_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n423_), .A3(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n459_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G71gat), .B(G99gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G43gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT31), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n457_), .B(KEYINPUT86), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n546_), .A3(new_n544_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n548_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n538_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n522_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n504_), .A2(new_n493_), .A3(new_n505_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(KEYINPUT100), .A3(new_n489_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT100), .B1(new_n559_), .B2(new_n489_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT27), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n445_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n379_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n567_));
  OAI22_X1  g366(.A1(new_n567_), .A2(KEYINPUT99), .B1(new_n434_), .B2(new_n509_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n568_), .B2(new_n519_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n564_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n556_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n554_), .A2(new_n555_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n537_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n535_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n563_), .A2(new_n565_), .A3(new_n571_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n558_), .A2(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n300_), .A2(new_n376_), .A3(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n563_), .A2(KEYINPUT101), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n559_), .A2(new_n489_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT100), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n560_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n579_), .A2(new_n272_), .A3(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n590_));
  AND2_X1   g389(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n376_), .A2(KEYINPUT102), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n571_), .A2(new_n565_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n576_), .A2(new_n583_), .A3(new_n560_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n595_), .A2(new_n596_), .B1(new_n522_), .B2(new_n557_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n262_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n376_), .A2(KEYINPUT102), .ZN(new_n600_));
  AND4_X1   g399(.A1(new_n593_), .A2(new_n599_), .A3(new_n600_), .A4(new_n298_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n584_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(G1gat), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n592_), .B(new_n603_), .C1(new_n590_), .C2(new_n589_), .ZN(G1324gat));
  NAND3_X1  g403(.A1(new_n579_), .A2(new_n273_), .A3(new_n594_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n594_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G8gat), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(G1325gat));
  NAND2_X1  g411(.A1(new_n601_), .A2(new_n556_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(G15gat), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT41), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n579_), .A2(new_n540_), .A3(new_n556_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT104), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(KEYINPUT41), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n617_), .A3(new_n618_), .ZN(G1326gat));
  INV_X1    g418(.A(G22gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n601_), .B2(new_n538_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT42), .Z(new_n622_));
  NAND3_X1  g421(.A1(new_n579_), .A2(new_n620_), .A3(new_n538_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1327gat));
  NAND4_X1  g423(.A1(new_n578_), .A2(new_n376_), .A3(new_n297_), .A4(new_n598_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n584_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n593_), .A2(new_n600_), .A3(new_n297_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT105), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  INV_X1    g430(.A(new_n263_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n576_), .A2(new_n583_), .A3(new_n560_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n594_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n557_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n446_), .A2(new_n447_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n636_), .A2(new_n500_), .A3(new_n499_), .A4(new_n491_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n568_), .A2(new_n519_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n581_), .B(new_n503_), .C1(new_n638_), .C2(new_n502_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n631_), .B(new_n632_), .C1(new_n634_), .C2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT43), .B1(new_n597_), .B2(new_n263_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n578_), .A2(KEYINPUT106), .A3(new_n631_), .A4(new_n632_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n628_), .B1(new_n630_), .B2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n629_), .A2(KEYINPUT105), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n629_), .A2(KEYINPUT105), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n646_), .B(KEYINPUT44), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n630_), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n646_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n588_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n627_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n654_), .B2(new_n594_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n594_), .A2(new_n658_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n625_), .A2(KEYINPUT109), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT109), .B1(new_n625_), .B2(new_n660_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n663_));
  AND3_X1   g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n657_), .B1(new_n659_), .B2(new_n667_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n595_), .B(new_n647_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n658_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1329gat));
  AOI21_X1  g470(.A(G43gat), .B1(new_n626_), .B2(new_n556_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n556_), .A2(G43gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n654_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1330gat));
  AOI21_X1  g475(.A(G50gat), .B1(new_n626_), .B2(new_n538_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n538_), .A2(G50gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n654_), .B2(new_n678_), .ZN(G1331gat));
  NAND2_X1  g478(.A1(new_n363_), .A2(new_n375_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AND4_X1   g480(.A1(new_n321_), .A2(new_n300_), .A3(new_n681_), .A4(new_n578_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n588_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n321_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n599_), .A2(new_n681_), .A3(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT111), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n584_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n689_), .B2(new_n683_), .ZN(G1332gat));
  INV_X1    g489(.A(G64gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n691_), .A3(new_n594_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n594_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G64gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT48), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT48), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n682_), .A2(new_n698_), .A3(new_n556_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n688_), .A2(new_n556_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G71gat), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n538_), .A2(new_n524_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT112), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n682_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n688_), .A2(new_n538_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G78gat), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n680_), .A2(new_n320_), .A3(new_n298_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n646_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n563_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n597_), .A2(new_n320_), .A3(new_n262_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n716_), .A2(new_n681_), .A3(new_n297_), .ZN(new_n717_));
  INV_X1    g516(.A(G85gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n588_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT113), .Z(G1336gat));
  AOI21_X1  g520(.A(G92gat), .B1(new_n717_), .B2(new_n594_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n714_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n594_), .A2(new_n227_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(G1337gat));
  AOI21_X1  g524(.A(new_n204_), .B1(new_n723_), .B2(new_n556_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n556_), .A2(new_n232_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n717_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1338gat));
  INV_X1    g529(.A(new_n538_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G106gat), .B1(new_n714_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n731_), .A2(G106gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n717_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n732_), .A2(new_n733_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g540(.A(KEYINPUT116), .B1(new_n680_), .B2(new_n686_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n743_), .B(new_n685_), .C1(new_n363_), .C2(new_n375_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n263_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(new_n263_), .C1(new_n742_), .C2(new_n744_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n318_), .A2(new_n319_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n327_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT117), .B1(new_n751_), .B2(new_n328_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n327_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n344_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n348_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n334_), .A2(KEYINPUT55), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n752_), .A2(new_n755_), .A3(new_n757_), .A4(new_n758_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n326_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n749_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT118), .B(new_n749_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n317_), .B1(new_n311_), .B2(new_n308_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n308_), .B2(new_n306_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n319_), .B(new_n767_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n765_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n262_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(KEYINPUT57), .A3(new_n262_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n761_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n759_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n326_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n359_), .A2(new_n319_), .A3(new_n767_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT120), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(KEYINPUT120), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n784_), .A3(new_n780_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n632_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n772_), .A2(new_n773_), .A3(new_n786_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n746_), .A2(new_n748_), .B1(new_n787_), .B2(new_n297_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n587_), .A2(new_n594_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n572_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n320_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n746_), .A2(new_n748_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n297_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n791_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT59), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT59), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n791_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(KEYINPUT59), .A3(new_n798_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT121), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n320_), .A2(G113gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT122), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n793_), .B1(new_n806_), .B2(new_n808_), .ZN(G1340gat));
  OR2_X1    g608(.A1(new_n680_), .A2(KEYINPUT60), .ZN(new_n810_));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n792_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n680_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n811_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT123), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n792_), .B2(new_n298_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n298_), .A2(G127gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT124), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n806_), .B2(new_n819_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n263_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n802_), .A2(new_n805_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n792_), .A2(new_n598_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n823_), .A2(KEYINPUT125), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1343gat));
  NOR2_X1   g629(.A1(new_n788_), .A2(new_n575_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n789_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n320_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n681_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g636(.A1(new_n832_), .A2(new_n297_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT61), .B(G155gat), .Z(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n832_), .B2(new_n263_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n262_), .A2(G162gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n832_), .B2(new_n842_), .ZN(G1347gat));
  NAND3_X1  g642(.A1(new_n587_), .A2(new_n594_), .A3(new_n790_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n788_), .A2(new_n321_), .A3(new_n399_), .A4(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n788_), .A2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n416_), .B1(new_n846_), .B2(new_n320_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(KEYINPUT62), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(KEYINPUT62), .B2(new_n847_), .ZN(G1348gat));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n681_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n298_), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n388_), .B(G183gat), .S(new_n852_), .Z(G1350gat));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n598_), .A3(new_n389_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n788_), .A2(new_n263_), .A3(new_n844_), .ZN(new_n855_));
  INV_X1    g654(.A(G190gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1351gat));
  NOR2_X1   g656(.A1(new_n595_), .A2(new_n584_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n831_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n321_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n402_), .ZN(G1352gat));
  INV_X1    g660(.A(new_n859_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n681_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n298_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n865_), .B2(new_n866_), .ZN(G1354gat));
  XOR2_X1   g668(.A(KEYINPUT126), .B(G218gat), .Z(new_n870_));
  NOR3_X1   g669(.A1(new_n859_), .A2(new_n263_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n862_), .A2(new_n598_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(G1355gat));
endmodule


