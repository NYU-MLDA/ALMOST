//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XOR2_X1   g002(.A(G211gat), .B(G218gat), .Z(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT90), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT89), .B(G204gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(new_n205_), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G197gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n204_), .B1(new_n215_), .B2(KEYINPUT21), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n213_), .B2(G197gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n206_), .A2(new_n207_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(G197gat), .ZN(new_n221_));
  NOR4_X1   g020(.A1(new_n206_), .A2(new_n207_), .A3(new_n218_), .A4(new_n205_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n217_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT92), .ZN(new_n224_));
  INV_X1    g023(.A(new_n207_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(KEYINPUT91), .A3(G197gat), .A4(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n206_), .A2(new_n207_), .A3(new_n205_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n219_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT92), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n217_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n216_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n204_), .A2(KEYINPUT21), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n238_));
  INV_X1    g037(.A(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI22_X1  g040(.A1(new_n237_), .A2(new_n238_), .B1(KEYINPUT24), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT82), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(G190gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT26), .B(G190gat), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(new_n243_), .ZN(new_n247_));
  OR2_X1    g046(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n242_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n241_), .A2(KEYINPUT24), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n255_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n256_), .B(KEYINPUT83), .ZN(new_n261_));
  INV_X1    g060(.A(new_n259_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT84), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n251_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n236_), .B(KEYINPUT23), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n258_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT85), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n239_), .B2(KEYINPUT22), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n240_), .B(new_n270_), .C1(new_n271_), .C2(new_n269_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n254_), .A2(new_n264_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n232_), .A2(new_n235_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT20), .ZN(new_n275_));
  AND2_X1   g074(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT97), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT97), .ZN(new_n279_));
  NAND2_X1  g078(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n248_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n246_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n259_), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT98), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n278_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n246_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT98), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n262_), .A2(new_n256_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n242_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n258_), .B1(new_n240_), .B2(new_n271_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n237_), .A2(new_n238_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n232_), .A2(new_n235_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n203_), .B1(new_n275_), .B2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G8gat), .B(G36gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n232_), .A2(new_n235_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n273_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n203_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n232_), .A2(new_n235_), .A3(new_n292_), .A4(new_n296_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n306_), .A2(KEYINPUT20), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n298_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n303_), .B1(new_n298_), .B2(new_n309_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n303_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n275_), .A2(new_n297_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n307_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n273_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(KEYINPUT20), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT104), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT20), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n292_), .A2(new_n296_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n219_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n210_), .B2(new_n205_), .ZN(new_n325_));
  AOI211_X1 g124(.A(KEYINPUT92), .B(KEYINPUT21), .C1(new_n325_), .C2(new_n227_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n230_), .B1(new_n229_), .B2(new_n217_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n234_), .B1(new_n328_), .B2(new_n216_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n322_), .B1(new_n323_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT104), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n307_), .B1(new_n321_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT105), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n317_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  AOI211_X1 g133(.A(KEYINPUT105), .B(new_n307_), .C1(new_n321_), .C2(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n315_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n298_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT27), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n314_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G155gat), .B(G162gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(G141gat), .ZN(new_n345_));
  INV_X1    g144(.A(G148gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT3), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT87), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n344_), .A2(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n351_), .A2(KEYINPUT87), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n342_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n346_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n342_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT88), .B1(new_n355_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n344_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n348_), .A2(new_n349_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n354_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n356_), .A2(new_n352_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n368_), .B(new_n357_), .C1(KEYINPUT1), .C2(new_n342_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n341_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n362_), .C2(new_n370_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G22gat), .B(G50gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n362_), .A2(new_n370_), .A3(KEYINPUT29), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n304_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n355_), .A2(new_n361_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n372_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n304_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT93), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT94), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n384_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(G228gat), .B(G233gat), .C1(new_n329_), .C2(new_n386_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n304_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n381_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n393_), .A2(new_n381_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(KEYINPUT95), .A3(new_n395_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n390_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n398_), .A2(new_n402_), .A3(KEYINPUT96), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT96), .B1(new_n398_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n397_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n340_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G113gat), .B(G120gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n408_), .A2(new_n409_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n362_), .A2(new_n370_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(KEYINPUT100), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT100), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n385_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n417_), .A3(KEYINPUT4), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n362_), .A2(new_n370_), .A3(new_n419_), .A4(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT101), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT102), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT102), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n418_), .A2(new_n426_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G85gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n424_), .A2(new_n434_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n273_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(G15gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(new_n412_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n442_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n407_), .A2(new_n436_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT103), .ZN(new_n450_));
  INV_X1    g249(.A(new_n309_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n322_), .B1(new_n329_), .B2(new_n273_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n297_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n307_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n315_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n432_), .A2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .A4(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n420_), .A2(new_n421_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n459_), .A2(new_n418_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n413_), .A2(new_n417_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n422_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n432_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n455_), .A2(new_n337_), .A3(new_n458_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n435_), .A2(new_n456_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n450_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n310_), .A2(new_n311_), .A3(new_n464_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT103), .A3(new_n467_), .A4(new_n458_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n472_));
  INV_X1    g271(.A(new_n317_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n306_), .B1(new_n330_), .B2(KEYINPUT104), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n319_), .A2(new_n320_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n203_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n473_), .B1(new_n476_), .B2(KEYINPUT105), .ZN(new_n477_));
  INV_X1    g276(.A(new_n335_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n472_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n298_), .A2(new_n309_), .A3(new_n472_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n436_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n469_), .B(new_n471_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n400_), .A2(new_n401_), .A3(new_n390_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n394_), .A2(new_n395_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n378_), .B(new_n380_), .C1(new_n485_), .C2(new_n392_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n483_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n398_), .A2(new_n402_), .A3(KEYINPUT96), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n436_), .B1(new_n489_), .B2(new_n397_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n482_), .A2(new_n406_), .B1(new_n490_), .B2(new_n340_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT107), .B1(new_n491_), .B2(new_n447_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT107), .ZN(new_n493_));
  INV_X1    g292(.A(new_n472_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n481_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n312_), .A2(new_n467_), .A3(new_n458_), .A4(new_n465_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n495_), .A2(new_n496_), .B1(new_n497_), .B2(new_n450_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n405_), .B1(new_n498_), .B2(new_n471_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n314_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n303_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n338_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n436_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n405_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n493_), .B(new_n448_), .C1(new_n499_), .C2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n449_), .B1(new_n492_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT65), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT66), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT6), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G85gat), .B(G92gat), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(KEYINPUT68), .A3(new_n520_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT8), .A3(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n519_), .A2(KEYINPUT67), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(KEYINPUT67), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n528_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT10), .B(G99gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n511_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n534_), .A2(new_n518_), .A3(new_n535_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G29gat), .B(G36gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G43gat), .B(G50gat), .Z(new_n544_));
  OR3_X1    g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT15), .Z(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  OAI221_X1 g350(.A(new_n549_), .B1(KEYINPUT35), .B2(new_n551_), .C1(new_n547_), .C2(new_n539_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT35), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT72), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n552_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n555_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n555_), .A2(new_n559_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n507_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT71), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT11), .Z(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT69), .B(G71gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G78gat), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(KEYINPUT11), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n539_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n531_), .A2(new_n575_), .A3(new_n577_), .A4(new_n538_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(KEYINPUT12), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n539_), .A2(new_n582_), .A3(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n580_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n570_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n589_), .A3(new_n570_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n547_), .B(KEYINPUT78), .ZN(new_n599_));
  INV_X1    g398(.A(G1gat), .ZN(new_n600_));
  INV_X1    g399(.A(G8gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT14), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n604_), .B(KEYINPUT14), .C1(new_n600_), .C2(new_n601_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G15gat), .B(G22gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT75), .ZN(new_n608_));
  XOR2_X1   g407(.A(G1gat), .B(G8gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n599_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT80), .ZN(new_n615_));
  INV_X1    g414(.A(new_n610_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n548_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n599_), .A2(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n612_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n614_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT79), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n615_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n620_), .A2(new_n626_), .B1(KEYINPUT79), .B2(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n598_), .A2(KEYINPUT111), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT111), .ZN(new_n632_));
  INV_X1    g431(.A(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n597_), .B2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n578_), .B(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n610_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT77), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT17), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n640_), .B(new_n646_), .Z(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(KEYINPUT17), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n638_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n564_), .A2(new_n635_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n503_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT112), .Z(new_n653_));
  NOR2_X1   g452(.A1(new_n507_), .A2(new_n633_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n563_), .B(KEYINPUT37), .ZN(new_n655_));
  INV_X1    g454(.A(new_n650_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n655_), .A2(new_n597_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT110), .B(KEYINPUT38), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n436_), .B(KEYINPUT109), .Z(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n600_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n653_), .A2(new_n663_), .A3(new_n664_), .ZN(G1324gat));
  OAI21_X1  g464(.A(G8gat), .B1(new_n651_), .B2(new_n340_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n502_), .A2(new_n601_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n667_), .A2(new_n668_), .B1(new_n659_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI221_X1 g471(.A(KEYINPUT40), .B1(new_n659_), .B2(new_n669_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n651_), .B2(new_n448_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n658_), .A2(G15gat), .A3(new_n448_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n406_), .A2(G22gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT113), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n654_), .A2(new_n657_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G22gat), .B1(new_n651_), .B2(new_n406_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(KEYINPUT42), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(KEYINPUT42), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT114), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT114), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n656_), .A2(new_n563_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT115), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n598_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n654_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n436_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n449_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n482_), .A2(new_n406_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n490_), .A2(new_n340_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n493_), .B1(new_n698_), .B2(new_n448_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n491_), .A2(KEYINPUT107), .A3(new_n447_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n655_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT37), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n563_), .B(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n507_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n631_), .A2(new_n656_), .A3(new_n634_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n711_), .B(new_n708_), .C1(new_n703_), .C2(new_n706_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n661_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n694_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n713_), .B2(new_n502_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n692_), .A2(new_n654_), .A3(new_n717_), .A4(new_n502_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n710_), .A2(new_n712_), .A3(new_n340_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT46), .B(new_n720_), .C1(new_n723_), .C2(new_n717_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1329gat));
  NOR4_X1   g524(.A1(new_n710_), .A2(new_n712_), .A3(new_n438_), .A4(new_n448_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G43gat), .B1(new_n693_), .B2(new_n447_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT47), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n448_), .A2(new_n438_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n713_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n693_), .B2(new_n405_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n405_), .A2(G50gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n713_), .B2(new_n735_), .ZN(G1331gat));
  NOR3_X1   g535(.A1(new_n598_), .A2(new_n630_), .A3(new_n656_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n564_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n503_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n701_), .A2(new_n633_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(KEYINPUT116), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n598_), .B1(new_n740_), .B2(KEYINPUT116), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n650_), .A3(new_n705_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n661_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(G57gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n744_), .B2(new_n746_), .ZN(G1332gat));
  OAI21_X1  g546(.A(G64gat), .B1(new_n738_), .B2(new_n340_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n340_), .A2(G64gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n744_), .B2(new_n750_), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n738_), .B2(new_n448_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n448_), .A2(G71gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n744_), .B2(new_n754_), .ZN(G1334gat));
  OR2_X1    g554(.A1(new_n406_), .A2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(G78gat), .B1(new_n738_), .B2(new_n406_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(KEYINPUT50), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(KEYINPUT50), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n744_), .A2(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(G1335gat));
  NAND3_X1  g559(.A1(new_n741_), .A2(new_n691_), .A3(new_n742_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G85gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n661_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n707_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n598_), .A2(new_n630_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n656_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n765_), .A2(new_n503_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n763_), .B2(new_n768_), .ZN(G1336gat));
  INV_X1    g568(.A(G92gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n762_), .A2(new_n770_), .A3(new_n502_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n765_), .A2(new_n340_), .A3(new_n767_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(new_n772_), .ZN(G1337gat));
  NOR2_X1   g572(.A1(new_n765_), .A2(new_n767_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n510_), .B1(new_n774_), .B2(new_n447_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n447_), .A2(new_n536_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n761_), .A2(new_n776_), .ZN(new_n777_));
  OR3_X1    g576(.A1(new_n775_), .A2(KEYINPUT51), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n775_), .B2(new_n777_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1338gat));
  NOR2_X1   g579(.A1(new_n406_), .A2(G106gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n743_), .A2(new_n691_), .A3(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n707_), .A2(new_n405_), .A3(new_n656_), .A4(new_n766_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(new_n782_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n586_), .A2(KEYINPUT117), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n584_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n581_), .A2(KEYINPUT118), .A3(new_n583_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n588_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n588_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT55), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n793_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n570_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT119), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n801_), .A2(new_n808_), .A3(KEYINPUT56), .A4(new_n802_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n592_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n624_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n611_), .A2(new_n612_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n617_), .A2(new_n618_), .A3(new_n613_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n614_), .A2(new_n619_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n814_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n810_), .B2(new_n590_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT120), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n593_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n813_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n563_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT57), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n563_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n819_), .A2(new_n592_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT58), .B1(new_n833_), .B2(KEYINPUT121), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n802_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n802_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n835_), .B(new_n836_), .C1(new_n839_), .C2(new_n832_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n840_), .A3(new_n655_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n828_), .A2(new_n831_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n656_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n705_), .A2(new_n598_), .A3(new_n633_), .A4(new_n650_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT54), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n407_), .A2(new_n745_), .A3(new_n448_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n630_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(KEYINPUT122), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n846_), .B(new_n847_), .C1(KEYINPUT122), .C2(KEYINPUT59), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n630_), .A2(G113gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT123), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n850_), .B1(new_n855_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n849_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n598_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n849_), .A2(new_n864_), .A3(new_n650_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n656_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n849_), .A2(new_n868_), .A3(new_n563_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n705_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1343gat));
  NOR3_X1   g670(.A1(new_n745_), .A2(new_n406_), .A3(new_n447_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n846_), .A2(new_n340_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n633_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n345_), .ZN(G1344gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n598_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n346_), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n873_), .A2(new_n656_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n873_), .B2(new_n705_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n827_), .A2(G162gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n873_), .B2(new_n882_), .ZN(G1347gat));
  NOR4_X1   g682(.A1(new_n340_), .A2(new_n661_), .A3(new_n405_), .A4(new_n448_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n846_), .A2(new_n630_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n239_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n885_), .B2(new_n239_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n271_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  AND2_X1   g689(.A1(new_n846_), .A2(new_n884_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n597_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n650_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n894_), .A2(new_n251_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n285_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n891_), .A2(new_n286_), .A3(new_n563_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n891_), .A2(new_n655_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n265_), .ZN(G1351gat));
  NAND2_X1  g699(.A1(new_n490_), .A2(new_n448_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(KEYINPUT124), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(KEYINPUT124), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n902_), .A2(new_n502_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(G197gat), .A3(new_n630_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n908_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G197gat), .B1(new_n906_), .B2(new_n630_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n906_), .A2(new_n597_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n220_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n213_), .B2(new_n913_), .ZN(G1353gat));
  AOI211_X1 g714(.A(KEYINPUT63), .B(G211gat), .C1(new_n906_), .C2(new_n650_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n846_), .A2(new_n904_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n917_), .A2(new_n656_), .A3(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n919_), .ZN(G1354gat));
  NAND2_X1  g719(.A1(new_n655_), .A2(G218gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT126), .Z(new_n922_));
  NOR2_X1   g721(.A1(new_n917_), .A2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G218gat), .B1(new_n906_), .B2(new_n563_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT127), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1355gat));
endmodule


