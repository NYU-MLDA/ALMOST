//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_;
  NAND2_X1  g000(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT25), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  OAI211_X1 g003(.A(KEYINPUT77), .B(G190gat), .C1(new_n204_), .C2(KEYINPUT76), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT76), .B1(new_n204_), .B2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT26), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .A4(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT78), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT24), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(new_n216_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(new_n214_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n214_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G227gat), .A2(G233gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT80), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G99gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n227_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G127gat), .B(G134gat), .Z(new_n233_));
  XOR2_X1   g032(.A(G113gat), .B(G120gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT79), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n236_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G1gat), .B(G29gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G85gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT3), .Z(new_n252_));
  NAND2_X1  g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT2), .Z(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n249_), .B1(new_n248_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n256_), .B2(new_n248_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n251_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n235_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n235_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n235_), .A2(new_n255_), .A3(KEYINPUT88), .A4(new_n260_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT4), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n247_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  AOI211_X1 g076(.A(new_n246_), .B(new_n275_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n242_), .A2(new_n279_), .ZN(new_n280_));
  OR3_X1    g079(.A1(new_n261_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT28), .B1(new_n261_), .B2(KEYINPUT29), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G22gat), .B(G50gat), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G204gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT82), .ZN(new_n294_));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295_));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n288_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n287_), .A2(KEYINPUT81), .A3(G197gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n290_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n295_), .B1(new_n299_), .B2(KEYINPUT21), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n291_), .B(KEYINPUT83), .Z(new_n301_));
  AND2_X1   g100(.A1(new_n295_), .A2(KEYINPUT21), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n294_), .A2(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n305_));
  OAI211_X1 g104(.A(G228gat), .B(G233gat), .C1(new_n303_), .C2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n294_), .A2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n302_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G78gat), .B(G106gat), .Z(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n286_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n314_), .B1(new_n316_), .B2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n306_), .A2(new_n312_), .A3(KEYINPUT84), .A4(new_n313_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n286_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AOI211_X1 g124(.A(KEYINPUT85), .B(new_n286_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n318_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT19), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n222_), .A2(KEYINPUT86), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT86), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n218_), .B(new_n334_), .C1(G183gat), .C2(G190gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n225_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G190gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n332_), .B1(new_n309_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n303_), .A2(new_n226_), .A3(new_n221_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n331_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  AND2_X1   g148(.A1(new_n336_), .A2(new_n340_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n332_), .B1(new_n350_), .B2(new_n303_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n309_), .A2(new_n227_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n331_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n345_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n349_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n351_), .A2(new_n331_), .A3(new_n352_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(new_n344_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n357_), .A3(KEYINPUT87), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT27), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n355_), .C1(new_n356_), .C2(new_n344_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n342_), .A2(new_n331_), .A3(new_n343_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n331_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n354_), .B(KEYINPUT27), .C1(new_n349_), .C2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n328_), .A2(new_n367_), .A3(KEYINPUT91), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT91), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n366_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n327_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n280_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n327_), .A2(new_n362_), .A3(new_n366_), .A4(new_n279_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT90), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n358_), .A2(new_n361_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n272_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n376_));
  AOI211_X1 g175(.A(new_n247_), .B(new_n376_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT33), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n274_), .A2(new_n247_), .A3(new_n276_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n278_), .A2(KEYINPUT33), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n277_), .A2(new_n278_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n365_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n345_), .A2(new_n353_), .A3(new_n384_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n365_), .B2(new_n384_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT89), .B1(new_n279_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n382_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n328_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n367_), .A2(new_n393_), .A3(new_n327_), .A4(new_n279_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n374_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n372_), .B1(new_n395_), .B2(new_n241_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G29gat), .B(G36gat), .Z(new_n397_));
  XOR2_X1   g196(.A(G43gat), .B(G50gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G22gat), .ZN(new_n401_));
  INV_X1    g200(.A(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(G8gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G8gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G229gat), .A2(G233gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n399_), .B(KEYINPUT15), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n407_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n400_), .B(new_n407_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n409_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n410_), .A2(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G113gat), .B(G141gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(G169gat), .B(G197gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n415_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n396_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G85gat), .ZN(new_n422_));
  INV_X1    g221(.A(G92gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT7), .ZN(new_n427_));
  INV_X1    g226(.A(G99gat), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT67), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n426_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n424_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n423_), .A2(KEYINPUT66), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G92gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n422_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT9), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT65), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT9), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n443_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n433_), .A2(new_n434_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT10), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT64), .B(G106gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G78gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT11), .ZN(new_n461_));
  XOR2_X1   g260(.A(G71gat), .B(G78gat), .Z(new_n462_));
  INV_X1    g261(.A(G64gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G57gat), .ZN(new_n464_));
  INV_X1    g263(.A(G57gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G64gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT11), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n461_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n424_), .A2(new_n471_), .A3(new_n425_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n436_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n440_), .A2(new_n458_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G230gat), .A2(G233gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n470_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n445_), .A2(G92gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n423_), .A2(KEYINPUT66), .ZN(new_n479_));
  OAI21_X1  g278(.A(G85gat), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n449_), .A2(new_n451_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n442_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n434_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT64), .B(G106gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n473_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n485_), .A2(KEYINPUT67), .A3(new_n435_), .A4(new_n430_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT8), .B1(new_n490_), .B2(new_n426_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n477_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT12), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n453_), .A2(new_n457_), .B1(new_n436_), .B2(new_n472_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n440_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n477_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n476_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n475_), .B1(new_n492_), .B2(new_n474_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G120gat), .B(G148gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G176gat), .B(G204gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n498_), .A2(new_n499_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT69), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(KEYINPUT13), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT70), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n515_), .A3(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n411_), .A2(new_n495_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n494_), .A2(new_n399_), .A3(new_n440_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT71), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n519_), .A2(new_n520_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(KEYINPUT71), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G134gat), .B(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT36), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n526_), .B(new_n527_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n531_), .B(KEYINPUT36), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT73), .ZN(new_n541_));
  XOR2_X1   g340(.A(G127gat), .B(G155gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT17), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n407_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n470_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(KEYINPUT17), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT74), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n539_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n421_), .A2(new_n518_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT38), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n383_), .A2(new_n402_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n537_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n396_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n518_), .A2(new_n567_), .A3(new_n419_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT93), .B1(new_n517_), .B2(new_n420_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n553_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(G1gat), .B1(new_n572_), .B2(new_n279_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n573_), .A3(new_n574_), .ZN(G1324gat));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n572_), .A2(new_n367_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n403_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT94), .B(G8gat), .C1(new_n572_), .C2(new_n367_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(KEYINPUT39), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n576_), .B(new_n581_), .C1(new_n577_), .C2(new_n403_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n559_), .A2(new_n403_), .A3(new_n370_), .A4(new_n560_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n580_), .A2(KEYINPUT40), .A3(new_n582_), .A4(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1325gat));
  OR2_X1    g387(.A1(new_n572_), .A2(new_n241_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G15gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT41), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(G15gat), .A3(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(KEYINPUT96), .A3(new_n594_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n241_), .A2(G15gat), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n561_), .A2(KEYINPUT97), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT97), .B1(new_n561_), .B2(new_n599_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .A4(new_n601_), .ZN(G1326gat));
  XOR2_X1   g401(.A(new_n327_), .B(KEYINPUT98), .Z(new_n603_));
  OAI21_X1  g402(.A(G22gat), .B1(new_n572_), .B2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT42), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n603_), .A2(G22gat), .ZN(new_n607_));
  OAI22_X1  g406(.A1(new_n605_), .A2(new_n606_), .B1(new_n561_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT99), .ZN(G1327gat));
  INV_X1    g408(.A(new_n539_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT43), .B1(new_n396_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT43), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n373_), .A2(KEYINPUT90), .B1(new_n391_), .B2(new_n328_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n242_), .B1(new_n613_), .B2(new_n394_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n612_), .B(new_n539_), .C1(new_n614_), .C2(new_n372_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n568_), .A2(new_n555_), .A3(new_n569_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT100), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(KEYINPUT44), .A3(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n383_), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(KEYINPUT101), .A3(G29gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT101), .B1(new_n623_), .B2(G29gat), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n421_), .A2(new_n518_), .A3(new_n555_), .A4(new_n565_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n279_), .A2(G29gat), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n625_), .A2(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n367_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(new_n622_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n370_), .B(KEYINPUT102), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(G36gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n627_), .A2(KEYINPUT45), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT45), .B1(new_n627_), .B2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(KEYINPUT46), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  INV_X1    g440(.A(new_n639_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n632_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1329gat));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n627_), .B2(new_n241_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n621_), .A2(G43gat), .A3(new_n242_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n622_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g449(.A(G50gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n627_), .B2(new_n603_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n621_), .A2(G50gat), .A3(new_n327_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n648_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT103), .ZN(G1331gat));
  NOR2_X1   g454(.A1(new_n396_), .A2(new_n419_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(new_n517_), .A3(new_n556_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n465_), .A3(new_n383_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n566_), .A2(new_n420_), .A3(new_n517_), .A4(new_n554_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n383_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n663_), .B2(new_n465_), .ZN(G1332gat));
  INV_X1    g463(.A(new_n634_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n463_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G64gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G64gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1333gat));
  INV_X1    g470(.A(G71gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n657_), .A2(new_n672_), .A3(new_n242_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n661_), .A2(new_n662_), .A3(new_n242_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT49), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G71gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G71gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1334gat));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n603_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n657_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n661_), .A2(new_n662_), .A3(new_n680_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(G78gat), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G78gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1335gat));
  NAND3_X1  g485(.A1(new_n555_), .A2(new_n517_), .A3(new_n420_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n611_), .B2(new_n615_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G85gat), .B1(new_n689_), .B2(new_n279_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n518_), .A2(new_n554_), .A3(new_n537_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n656_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n422_), .A3(new_n383_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1336gat));
  AOI21_X1  g494(.A(G92gat), .B1(new_n693_), .B2(new_n370_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n634_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n688_), .B2(new_n697_), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n689_), .B2(new_n241_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n241_), .A2(new_n487_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n693_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n701_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n692_), .A2(KEYINPUT106), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT107), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n705_), .B(new_n707_), .ZN(G1338gat));
  AOI21_X1  g507(.A(new_n429_), .B1(new_n688_), .B2(new_n327_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT110), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n328_), .B(new_n687_), .C1(new_n611_), .C2(new_n615_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n429_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n710_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n711_), .B(new_n714_), .C1(new_n712_), .C2(new_n429_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n328_), .A2(new_n486_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n692_), .A2(KEYINPUT108), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT108), .B1(new_n692_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT53), .B1(new_n716_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n710_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n725_), .A2(new_n717_), .A3(new_n726_), .A4(new_n722_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1339gat));
  NAND3_X1  g527(.A1(new_n554_), .A2(new_n420_), .A3(new_n513_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(KEYINPUT111), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT54), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n539_), .B1(new_n729_), .B2(KEYINPUT111), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n412_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n418_), .B1(new_n413_), .B2(new_n409_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n415_), .A2(new_n418_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n508_), .A2(KEYINPUT115), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT115), .B1(new_n508_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n419_), .A2(new_n506_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n474_), .A2(new_n475_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n496_), .B1(new_n495_), .B2(new_n477_), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT12), .B(new_n470_), .C1(new_n494_), .C2(new_n440_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n747_), .B(KEYINPUT55), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n474_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n475_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT112), .B1(new_n498_), .B2(KEYINPUT55), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n754_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n505_), .B1(new_n759_), .B2(KEYINPUT113), .ZN(new_n760_));
  INV_X1    g559(.A(new_n475_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n474_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n761_), .A2(new_n762_), .B1(new_n498_), .B2(KEYINPUT55), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n498_), .A2(KEYINPUT112), .A3(KEYINPUT55), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n760_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n504_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n759_), .A2(KEYINPUT113), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n746_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n744_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n769_), .B1(new_n760_), .B2(new_n768_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n772_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n745_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n565_), .B1(new_n776_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n737_), .B1(new_n781_), .B2(KEYINPUT57), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n740_), .A2(new_n506_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n539_), .B1(new_n784_), .B2(KEYINPUT58), .ZN(new_n785_));
  INV_X1    g584(.A(new_n783_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n781_), .B2(KEYINPUT57), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n743_), .B1(new_n779_), .B2(KEYINPUT114), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n775_), .B(new_n745_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n537_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT116), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n782_), .A2(new_n791_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n553_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n736_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n368_), .A2(new_n371_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n383_), .A3(new_n242_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n781_), .A2(KEYINPUT57), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT57), .B(new_n537_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n787_), .A2(new_n788_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n784_), .A2(KEYINPUT58), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n539_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n555_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n736_), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n801_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n803_), .A2(new_n419_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G113gat), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n420_), .A2(G113gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n802_), .B2(new_n819_), .ZN(G1340gat));
  NAND3_X1  g619(.A1(new_n803_), .A2(new_n517_), .A3(new_n816_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n518_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(KEYINPUT60), .B2(new_n823_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n822_), .B1(new_n802_), .B2(new_n825_), .ZN(G1341gat));
  NOR2_X1   g625(.A1(new_n799_), .A2(new_n801_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G127gat), .B1(new_n827_), .B2(new_n554_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n803_), .A2(new_n816_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n553_), .A2(G127gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT119), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n827_), .B2(new_n565_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT121), .B(G134gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n539_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT122), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n834_), .A2(new_n835_), .B1(new_n829_), .B2(new_n838_), .ZN(G1343gat));
  NAND3_X1  g638(.A1(new_n327_), .A2(new_n383_), .A3(new_n241_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n799_), .A2(new_n665_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n419_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n517_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n554_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n841_), .A2(new_n849_), .A3(new_n565_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n841_), .A2(new_n539_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1347gat));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  INV_X1    g652(.A(new_n280_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n665_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n680_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n813_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n420_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n858_), .B2(new_n213_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT62), .B(G169gat), .C1(new_n857_), .C2(new_n420_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n224_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(G1348gat));
  NOR3_X1   g661(.A1(new_n855_), .A2(new_n214_), .A3(new_n518_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n736_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n794_), .A2(KEYINPUT116), .A3(new_n795_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT116), .B1(new_n794_), .B2(new_n795_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n809_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n867_), .B2(new_n553_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT123), .B1(new_n868_), .B2(new_n328_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n799_), .A2(new_n870_), .A3(new_n327_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n863_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT124), .B(new_n863_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n813_), .A2(new_n517_), .A3(new_n856_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n214_), .B2(new_n876_), .ZN(G1349gat));
  NOR3_X1   g676(.A1(new_n857_), .A2(new_n338_), .A3(new_n798_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n665_), .A2(new_n854_), .A3(new_n554_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  AOI21_X1  g681(.A(G183gat), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT125), .B(new_n880_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n878_), .B1(new_n883_), .B2(new_n884_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n857_), .B2(new_n610_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n565_), .A2(new_n337_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n857_), .B2(new_n887_), .ZN(G1351gat));
  NAND3_X1  g687(.A1(new_n327_), .A2(new_n279_), .A3(new_n241_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n889_), .A2(KEYINPUT126), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(KEYINPUT126), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n799_), .A2(new_n634_), .A3(new_n890_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n419_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n517_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n895_), .B(new_n896_), .Z(G1353gat));
  NAND2_X1  g696(.A1(new_n892_), .A2(new_n553_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT63), .B(G211gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n898_), .B2(new_n901_), .ZN(G1354gat));
  INV_X1    g701(.A(G218gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n892_), .A2(new_n903_), .A3(new_n565_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n892_), .A2(new_n539_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1355gat));
endmodule


