//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1020_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1032_, new_n1033_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT0), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT99), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G57gat), .B(G85gat), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT90), .ZN(new_n214_));
  INV_X1    g013(.A(G155gat), .ZN(new_n215_));
  INV_X1    g014(.A(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT91), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n225_), .A3(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228_));
  INV_X1    g027(.A(G141gat), .ZN(new_n229_));
  INV_X1    g028(.A(G148gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n220_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n230_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n221_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n217_), .A2(new_n218_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n219_), .B(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n213_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT89), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n243_), .A2(new_n244_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n220_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n221_), .A2(new_n225_), .A3(new_n222_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n225_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n219_), .B(KEYINPUT1), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n217_), .A2(new_n218_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n221_), .B(new_n236_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n259_), .A3(KEYINPUT92), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(new_n250_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n249_), .A2(new_n245_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n261_), .A2(KEYINPUT4), .A3(new_n263_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n267_));
  NAND4_X1  g066(.A1(new_n242_), .A2(new_n260_), .A3(new_n250_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n264_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n212_), .B(new_n265_), .C1(new_n266_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT101), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(new_n263_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n269_), .B(new_n268_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT101), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n265_), .A4(new_n212_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n265_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n212_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT25), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G183gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT95), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n291_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(G190gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT26), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(KEYINPUT26), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(G190gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT96), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n292_), .A2(new_n295_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT23), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(G183gat), .A3(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT97), .B1(new_n305_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n292_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT95), .B1(new_n289_), .B2(new_n291_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT96), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT96), .B1(new_n302_), .B2(new_n303_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n321_), .A2(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT97), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n310_), .B1(G183gat), .B2(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n311_), .A2(KEYINPUT22), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G169gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n332_), .A3(new_n312_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n314_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n320_), .A2(new_n328_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT93), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(G197gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n337_), .A2(G197gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n339_), .A2(G204gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT21), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G218gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G211gat), .ZN(new_n348_));
  INV_X1    g147(.A(G211gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G218gat), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n341_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n287_), .B1(new_n335_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT94), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT94), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n307_), .A2(new_n309_), .B1(new_n317_), .B2(new_n316_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n302_), .A2(KEYINPUT87), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n289_), .A2(KEYINPUT85), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n299_), .A3(KEYINPUT26), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .A4(new_n303_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n291_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n290_), .A2(KEYINPUT86), .A3(G183gat), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n369_), .B(new_n370_), .C1(KEYINPUT85), .C2(new_n289_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n315_), .B(new_n362_), .C1(new_n367_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n333_), .A2(KEYINPUT88), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT88), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n330_), .A2(new_n332_), .A3(new_n374_), .A4(new_n312_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n329_), .A2(new_n314_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n361_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n286_), .B1(new_n357_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n352_), .A2(KEYINPUT94), .A3(new_n355_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT94), .B1(new_n352_), .B2(new_n355_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n356_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n320_), .A2(new_n385_), .A3(new_n328_), .A4(new_n334_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n285_), .A2(new_n287_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n379_), .A2(new_n389_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n328_), .A2(new_n334_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n326_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n356_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT20), .A3(new_n378_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n285_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n395_), .B1(new_n400_), .B2(new_n388_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n283_), .B1(new_n394_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT102), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n393_), .B1(new_n379_), .B2(new_n389_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n395_), .A3(new_n388_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT102), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n283_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n384_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n334_), .B1(new_n305_), .B2(new_n319_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT20), .B1(new_n410_), .B2(new_n356_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n285_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n399_), .B2(new_n285_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n393_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n394_), .A2(new_n283_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n403_), .A2(new_n408_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418_));
  INV_X1    g217(.A(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n420_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n417_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT31), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n426_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n250_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n428_), .A3(new_n250_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n242_), .A2(new_n260_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n436_), .A2(KEYINPUT28), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(KEYINPUT28), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G22gat), .B(G50gat), .Z(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n435_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n442_));
  OAI211_X1 g241(.A(G228gat), .B(G233gat), .C1(new_n442_), .C2(new_n385_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n242_), .A2(KEYINPUT29), .A3(new_n260_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G228gat), .A2(G233gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n359_), .A2(new_n447_), .A3(new_n360_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n443_), .B(new_n445_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n242_), .A2(KEYINPUT29), .A3(new_n260_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n447_), .A3(new_n382_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n445_), .B1(new_n452_), .B2(new_n443_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n441_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n443_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n449_), .A3(new_n440_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n439_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n439_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND4_X1   g260(.A1(new_n282_), .A2(new_n416_), .A3(new_n433_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n415_), .A2(new_n414_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n407_), .B1(new_n406_), .B2(new_n283_), .ZN(new_n464_));
  AOI211_X1 g263(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n404_), .C2(new_n405_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n282_), .A3(new_n460_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT103), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n403_), .A2(new_n408_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT103), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n454_), .A2(new_n439_), .A3(new_n457_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n471_), .A2(new_n458_), .A3(new_n281_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n470_), .A3(new_n472_), .A4(new_n463_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n413_), .A2(KEYINPUT32), .A3(new_n395_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n400_), .A2(new_n388_), .A3(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n281_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT100), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n271_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n273_), .A2(new_n269_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(new_n268_), .C1(new_n274_), .C2(new_n265_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n279_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n480_), .A2(new_n483_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n479_), .B1(new_n271_), .B2(new_n478_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n461_), .B1(new_n477_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n468_), .A2(new_n473_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n433_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n462_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G22gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G15gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n422_), .A2(G22gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT78), .ZN(new_n499_));
  XOR2_X1   g298(.A(G1gat), .B(G8gat), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n498_), .A2(KEYINPUT78), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(KEYINPUT78), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT82), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512_));
  AOI211_X1 g311(.A(new_n512_), .B(new_n509_), .C1(new_n502_), .C2(new_n505_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n502_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT81), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n502_), .A2(new_n517_), .A3(new_n505_), .A4(new_n509_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n491_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n506_), .A2(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n519_), .A2(new_n491_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT83), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n491_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n505_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n500_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n510_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n512_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n506_), .A2(KEYINPUT82), .A3(new_n510_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n516_), .A2(new_n518_), .B1(new_n506_), .B2(new_n521_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n491_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n524_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n520_), .A2(new_n523_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT84), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n524_), .B2(new_n537_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  XOR2_X1   g352(.A(G120gat), .B(G148gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  XOR2_X1   g357(.A(G85gat), .B(G92gat), .Z(new_n559_));
  INV_X1    g358(.A(KEYINPUT64), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(KEYINPUT9), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT10), .B(G99gat), .Z(new_n562_));
  INV_X1    g361(.A(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G85gat), .B1(KEYINPUT64), .B2(G92gat), .ZN(new_n565_));
  INV_X1    g364(.A(G92gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n561_), .A2(new_n564_), .A3(new_n569_), .A4(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT65), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT65), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT7), .ZN(new_n581_));
  INV_X1    g380(.A(G99gat), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .A4(new_n563_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n578_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT66), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n574_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(KEYINPUT66), .A3(new_n573_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n559_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT8), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT8), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n559_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n585_), .B2(new_n575_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n577_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT11), .ZN(new_n598_));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n597_), .A2(KEYINPUT11), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n596_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n592_), .B1(new_n589_), .B2(new_n559_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n576_), .B1(new_n607_), .B2(new_n594_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n604_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT12), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(KEYINPUT12), .A3(new_n604_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(new_n611_), .A3(new_n606_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(new_n617_), .A3(KEYINPUT67), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT67), .B1(new_n613_), .B2(new_n617_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT69), .B(new_n558_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n558_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT70), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT70), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n613_), .A2(new_n617_), .A3(new_n625_), .A4(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n620_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n618_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT69), .B1(new_n630_), .B2(new_n558_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n553_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n558_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT69), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(KEYINPUT13), .A3(new_n621_), .A4(new_n627_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n490_), .A2(new_n552_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n596_), .A2(new_n509_), .B1(new_n642_), .B2(new_n641_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT73), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n608_), .A2(new_n646_), .A3(new_n521_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n608_), .B2(new_n521_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(KEYINPUT72), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT72), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n608_), .A2(new_n521_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT73), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n647_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n652_), .B1(new_n655_), .B2(new_n645_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n644_), .B1(new_n651_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G190gat), .B(G218gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT74), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT36), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n650_), .A2(KEYINPUT72), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n655_), .A2(new_n652_), .A3(new_n645_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n643_), .A3(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n657_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n662_), .B(KEYINPUT36), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT75), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n657_), .B2(new_n667_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n668_), .A2(new_n671_), .A3(KEYINPUT105), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT75), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n669_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n667_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n643_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n657_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n673_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n672_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n506_), .B(new_n682_), .Z(new_n683_));
  INV_X1    g482(.A(KEYINPUT17), .ZN(new_n684_));
  XNOR2_X1  g483(.A(G127gat), .B(G155gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT16), .ZN(new_n686_));
  XNOR2_X1  g485(.A(G183gat), .B(G211gat), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n686_), .B(new_n687_), .Z(new_n688_));
  AOI22_X1  g487(.A1(new_n683_), .A2(new_n605_), .B1(new_n684_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n605_), .B2(new_n683_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n688_), .A2(KEYINPUT79), .A3(new_n684_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n690_), .B(new_n691_), .Z(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n681_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n638_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G1gat), .B1(new_n695_), .B2(new_n282_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n632_), .A2(KEYINPUT71), .A3(new_n636_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT71), .B1(new_n632_), .B2(new_n636_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT37), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT76), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n670_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n675_), .A2(KEYINPUT76), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n700_), .B1(new_n705_), .B2(new_n679_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n668_), .A2(new_n671_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n706_), .A2(KEYINPUT77), .B1(new_n707_), .B2(new_n700_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n706_), .A2(KEYINPUT77), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n693_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n699_), .A2(KEYINPUT80), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT80), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n697_), .A2(new_n698_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n706_), .A2(KEYINPUT77), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n707_), .A2(new_n700_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n706_), .A2(KEYINPUT77), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n692_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n712_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n490_), .A2(new_n552_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n711_), .A2(new_n719_), .A3(new_n720_), .A4(KEYINPUT104), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n723_), .A2(new_n492_), .A3(new_n281_), .A4(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT38), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT38), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n696_), .B1(new_n726_), .B2(new_n727_), .ZN(G1324gat));
  NAND4_X1  g527(.A1(new_n723_), .A2(new_n493_), .A3(new_n466_), .A4(new_n724_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT39), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(G8gat), .C1(new_n695_), .C2(new_n416_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n473_), .A2(new_n487_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n470_), .B1(new_n416_), .B2(new_n472_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n489_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n462_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n637_), .A2(new_n552_), .ZN(new_n737_));
  AND4_X1   g536(.A1(new_n694_), .A2(new_n736_), .A3(new_n466_), .A4(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT39), .B1(new_n738_), .B2(new_n493_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n731_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n729_), .A2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n742_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n740_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1325gat));
  INV_X1    g545(.A(new_n695_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n422_), .B1(new_n747_), .B2(new_n433_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT41), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n489_), .A2(G15gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n723_), .A2(new_n724_), .A3(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT107), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT107), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n750_), .B(new_n751_), .C1(new_n754_), .C2(new_n755_), .ZN(G1326gat));
  OAI21_X1  g555(.A(G22gat), .B1(new_n695_), .B2(new_n461_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n461_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n723_), .A2(new_n495_), .A3(new_n760_), .A4(new_n724_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1327gat));
  NOR2_X1   g561(.A1(new_n672_), .A2(new_n680_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n692_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n638_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G29gat), .B1(new_n766_), .B2(new_n281_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n737_), .A2(new_n693_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n716_), .A2(new_n717_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n736_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n708_), .A2(new_n709_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n490_), .A2(new_n773_), .A3(KEYINPUT43), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n777_), .A2(G29gat), .A3(new_n281_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n736_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n773_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n768_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT44), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n767_), .B1(new_n778_), .B2(new_n782_), .ZN(G1328gat));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n784_));
  INV_X1    g583(.A(G36gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n416_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n782_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n638_), .A2(new_n785_), .A3(new_n466_), .A4(new_n764_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n784_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n466_), .B1(new_n781_), .B2(KEYINPUT44), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n775_), .A2(new_n776_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G36gat), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n788_), .B(new_n789_), .Z(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(KEYINPUT46), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n796_), .ZN(G1329gat));
  NAND4_X1  g596(.A1(new_n777_), .A2(new_n782_), .A3(G43gat), .A4(new_n433_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n419_), .B1(new_n765_), .B2(new_n489_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1330gat));
  NOR2_X1   g602(.A1(new_n461_), .A2(G50gat), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT112), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n766_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n777_), .A2(new_n760_), .A3(new_n782_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT111), .B1(new_n807_), .B2(G50gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n808_), .B2(new_n809_), .ZN(G1331gat));
  INV_X1    g609(.A(new_n637_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n718_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n551_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n710_), .A2(new_n814_), .A3(new_n637_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n812_), .A2(KEYINPUT114), .A3(new_n815_), .A4(new_n813_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(G57gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n281_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n813_), .A2(new_n713_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n694_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G57gat), .B1(new_n824_), .B2(new_n282_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1332gat));
  INV_X1    g625(.A(G64gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n827_), .A3(new_n466_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT48), .ZN(new_n829_));
  INV_X1    g628(.A(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n466_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(G64gat), .ZN(new_n832_));
  AOI211_X1 g631(.A(KEYINPUT48), .B(new_n827_), .C1(new_n830_), .C2(new_n466_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n832_), .B2(new_n833_), .ZN(G1333gat));
  XOR2_X1   g633(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n835_));
  NAND4_X1  g634(.A1(new_n813_), .A2(new_n694_), .A3(new_n433_), .A4(new_n713_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(G71gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n836_), .B2(G71gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(G71gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT116), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n836_), .A2(new_n837_), .A3(G71gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n835_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n489_), .A2(G71gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n818_), .A2(new_n819_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT117), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n840_), .A2(new_n845_), .A3(new_n847_), .A4(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1334gat));
  INV_X1    g651(.A(G78gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n820_), .A2(new_n853_), .A3(new_n760_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G78gat), .B1(new_n824_), .B2(new_n461_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n856_));
  OR2_X1    g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n856_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n857_), .A3(new_n858_), .ZN(G1335gat));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n551_), .A2(new_n692_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n637_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n637_), .B2(new_n861_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G85gat), .B1(new_n865_), .B2(new_n282_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n823_), .A2(new_n764_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n282_), .A2(G85gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1336gat));
  OAI21_X1  g668(.A(G92gat), .B1(new_n865_), .B2(new_n416_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n466_), .A2(new_n566_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n867_), .B2(new_n871_), .ZN(G1337gat));
  INV_X1    g671(.A(new_n865_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n582_), .B1(new_n873_), .B2(new_n433_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n562_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n867_), .A2(new_n875_), .A3(new_n489_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT120), .B(KEYINPUT51), .Z(new_n877_));
  OR3_X1    g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1338gat));
  NAND4_X1  g679(.A1(new_n823_), .A2(new_n563_), .A3(new_n760_), .A4(new_n764_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n760_), .B(new_n864_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n882_), .A2(new_n883_), .A3(G106gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(G106gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n881_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT53), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n881_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1339gat));
  NAND2_X1  g689(.A1(new_n811_), .A2(new_n552_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n718_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n710_), .A2(new_n893_), .A3(new_n552_), .A4(new_n811_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n547_), .A2(new_n550_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n617_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT55), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n617_), .A2(new_n898_), .A3(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n615_), .A2(new_n606_), .A3(new_n616_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n612_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n902_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n558_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n635_), .A2(new_n621_), .A3(new_n627_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n491_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n544_), .B1(new_n535_), .B2(new_n525_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n543_), .A2(new_n544_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n897_), .A2(new_n910_), .B1(new_n911_), .B2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n896_), .B1(new_n915_), .B2(new_n681_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n627_), .A2(new_n914_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n910_), .B2(new_n919_), .ZN(new_n920_));
  AOI211_X1 g719(.A(KEYINPUT58), .B(new_n918_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n709_), .B(new_n708_), .C1(new_n920_), .C2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n914_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n909_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n905_), .B2(new_n558_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n548_), .A2(new_n545_), .ZN(new_n927_));
  AOI211_X1 g726(.A(KEYINPUT84), .B(new_n544_), .C1(new_n524_), .C2(new_n537_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n627_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n923_), .B1(new_n926_), .B2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n930_), .A2(KEYINPUT57), .A3(new_n763_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n916_), .A2(new_n922_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n693_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n895_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n935_));
  NOR4_X1   g734(.A1(new_n489_), .A2(new_n466_), .A3(new_n760_), .A4(new_n282_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  AOI21_X1  g737(.A(KEYINPUT57), .B1(new_n930_), .B2(new_n763_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n922_), .B(new_n931_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n916_), .A2(KEYINPUT122), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n693_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n938_), .B1(new_n943_), .B2(new_n895_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n937_), .B1(new_n944_), .B2(new_n935_), .ZN(new_n945_));
  OAI21_X1  g744(.A(G113gat), .B1(new_n945_), .B2(new_n552_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n895_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n936_), .ZN(new_n948_));
  OR3_X1    g747(.A1(new_n948_), .A2(G113gat), .A3(new_n552_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1340gat));
  OAI21_X1  g749(.A(G120gat), .B1(new_n945_), .B2(new_n699_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n811_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n944_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n954_), .ZN(G1341gat));
  OAI21_X1  g754(.A(G127gat), .B1(new_n945_), .B2(new_n693_), .ZN(new_n956_));
  OR3_X1    g755(.A1(new_n948_), .A2(G127gat), .A3(new_n693_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1342gat));
  OAI21_X1  g757(.A(G134gat), .B1(new_n945_), .B2(new_n773_), .ZN(new_n959_));
  OR3_X1    g758(.A1(new_n948_), .A2(G134gat), .A3(new_n763_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1343gat));
  NAND3_X1  g760(.A1(new_n489_), .A2(new_n281_), .A3(new_n760_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n466_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n964_), .B1(new_n943_), .B2(new_n895_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n551_), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT123), .B(G141gat), .Z(new_n967_));
  XNOR2_X1  g766(.A(new_n966_), .B(new_n967_), .ZN(G1344gat));
  NAND2_X1  g767(.A1(new_n965_), .A2(new_n713_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g769(.A1(new_n965_), .A2(new_n692_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(KEYINPUT61), .B(G155gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1346gat));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n216_), .B1(new_n965_), .B2(new_n771_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n681_), .A2(new_n216_), .ZN(new_n976_));
  AOI211_X1 g775(.A(new_n964_), .B(new_n976_), .C1(new_n943_), .C2(new_n895_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n974_), .B1(new_n975_), .B2(new_n977_), .ZN(new_n978_));
  NAND4_X1  g777(.A1(new_n947_), .A2(new_n216_), .A3(new_n681_), .A4(new_n963_), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n773_), .B(new_n964_), .C1(new_n943_), .C2(new_n895_), .ZN(new_n980_));
  OAI211_X1 g779(.A(new_n979_), .B(KEYINPUT124), .C1(new_n980_), .C2(new_n216_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n978_), .A2(new_n981_), .ZN(G1347gat));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n489_), .A2(new_n281_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n466_), .ZN(new_n985_));
  INV_X1    g784(.A(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(new_n461_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n987_), .B1(new_n895_), .B2(new_n933_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n988_), .A2(new_n551_), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n983_), .B1(new_n989_), .B2(G169gat), .ZN(new_n990_));
  AOI211_X1 g789(.A(KEYINPUT62), .B(new_n311_), .C1(new_n988_), .C2(new_n551_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n330_), .A2(new_n332_), .ZN(new_n992_));
  OAI22_X1  g791(.A1(new_n990_), .A2(new_n991_), .B1(new_n992_), .B2(new_n989_), .ZN(G1348gat));
  AOI21_X1  g792(.A(G176gat), .B1(new_n988_), .B2(new_n637_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n947_), .A2(new_n461_), .ZN(new_n995_));
  INV_X1    g794(.A(new_n995_), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n699_), .A2(new_n312_), .A3(new_n985_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n994_), .B1(new_n996_), .B2(new_n997_), .ZN(G1349gat));
  NAND2_X1  g797(.A1(new_n986_), .A2(new_n692_), .ZN(new_n999_));
  AOI211_X1 g798(.A(new_n760_), .B(new_n999_), .C1(new_n943_), .C2(new_n895_), .ZN(new_n1000_));
  AOI21_X1  g799(.A(G183gat), .B1(new_n1000_), .B2(KEYINPUT125), .ZN(new_n1001_));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1002_), .B1(new_n995_), .B2(new_n999_), .ZN(new_n1003_));
  NOR3_X1   g802(.A1(new_n693_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n1004_));
  AOI22_X1  g803(.A1(new_n1001_), .A2(new_n1003_), .B1(new_n988_), .B2(new_n1004_), .ZN(G1350gat));
  NAND2_X1  g804(.A1(new_n301_), .A2(new_n304_), .ZN(new_n1006_));
  NAND3_X1  g805(.A1(new_n988_), .A2(new_n681_), .A3(new_n1006_), .ZN(new_n1007_));
  INV_X1    g806(.A(new_n1007_), .ZN(new_n1008_));
  AOI21_X1  g807(.A(new_n299_), .B1(new_n988_), .B2(new_n771_), .ZN(new_n1009_));
  OAI21_X1  g808(.A(KEYINPUT126), .B1(new_n1008_), .B2(new_n1009_), .ZN(new_n1010_));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n1011_));
  AND2_X1   g810(.A1(new_n988_), .A2(new_n771_), .ZN(new_n1012_));
  OAI211_X1 g811(.A(new_n1007_), .B(new_n1011_), .C1(new_n1012_), .C2(new_n299_), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(new_n1010_), .A2(new_n1013_), .ZN(G1351gat));
  NOR3_X1   g813(.A1(new_n416_), .A2(new_n433_), .A3(new_n467_), .ZN(new_n1015_));
  INV_X1    g814(.A(new_n1015_), .ZN(new_n1016_));
  AOI21_X1  g815(.A(new_n1016_), .B1(new_n943_), .B2(new_n895_), .ZN(new_n1017_));
  NAND2_X1  g816(.A1(new_n1017_), .A2(new_n551_), .ZN(new_n1018_));
  XNOR2_X1  g817(.A(new_n1018_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g818(.A1(new_n1017_), .A2(new_n713_), .ZN(new_n1020_));
  XNOR2_X1  g819(.A(new_n1020_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g820(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1022_));
  INV_X1    g821(.A(new_n1022_), .ZN(new_n1023_));
  NAND2_X1  g822(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1024_));
  AND4_X1   g823(.A1(new_n692_), .A2(new_n1017_), .A3(new_n1023_), .A4(new_n1024_), .ZN(new_n1025_));
  AOI211_X1 g824(.A(new_n693_), .B(new_n1016_), .C1(new_n943_), .C2(new_n895_), .ZN(new_n1026_));
  OAI21_X1  g825(.A(KEYINPUT127), .B1(new_n1026_), .B2(new_n1023_), .ZN(new_n1027_));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1028_));
  NAND2_X1  g827(.A1(new_n947_), .A2(new_n1015_), .ZN(new_n1029_));
  OAI211_X1 g828(.A(new_n1028_), .B(new_n1022_), .C1(new_n1029_), .C2(new_n693_), .ZN(new_n1030_));
  AOI21_X1  g829(.A(new_n1025_), .B1(new_n1027_), .B2(new_n1030_), .ZN(G1354gat));
  OAI21_X1  g830(.A(G218gat), .B1(new_n1029_), .B2(new_n773_), .ZN(new_n1032_));
  NAND3_X1  g831(.A1(new_n1017_), .A2(new_n347_), .A3(new_n681_), .ZN(new_n1033_));
  NAND2_X1  g832(.A1(new_n1032_), .A2(new_n1033_), .ZN(G1355gat));
endmodule


