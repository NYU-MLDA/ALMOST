//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT84), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT84), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(G155gat), .ZN(new_n211_));
  INV_X1    g010(.A(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n203_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n205_), .A2(new_n207_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n215_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n202_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n202_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n231_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G78gat), .B(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT88), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243_));
  INV_X1    g042(.A(G211gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G218gat), .ZN(new_n245_));
  INV_X1    g044(.A(G218gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G211gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(G211gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(G218gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT87), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT86), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G197gat), .B(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n254_), .A2(new_n255_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n262_), .A2(KEYINPUT85), .B1(G228gat), .B2(G233gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n262_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n234_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n242_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n242_), .B2(new_n267_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271_));
  INV_X1    g070(.A(G183gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT25), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G183gat), .ZN(new_n275_));
  INV_X1    g074(.A(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT26), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT26), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G190gat), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n273_), .A2(new_n275_), .A3(new_n277_), .A4(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT89), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291_));
  INV_X1    g090(.A(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n286_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n298_), .A3(new_n287_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT89), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n285_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n272_), .A2(new_n276_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n287_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT90), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n298_), .A2(new_n302_), .A3(KEYINPUT90), .A4(new_n287_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n260_), .A2(new_n301_), .A3(new_n261_), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n303_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n280_), .A2(new_n284_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n299_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n252_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n258_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n316_), .A3(KEYINPUT20), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n290_), .A2(new_n286_), .A3(new_n294_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n299_), .A2(KEYINPUT89), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n312_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n325_));
  OAI22_X1  g124(.A1(new_n314_), .A2(new_n315_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n312_), .A2(new_n299_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n260_), .A2(new_n261_), .A3(new_n327_), .A4(new_n311_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT20), .A4(new_n319_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n271_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT95), .B1(new_n324_), .B2(new_n325_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT95), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n301_), .A2(new_n338_), .A3(new_n309_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n314_), .A2(new_n315_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT96), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT20), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n316_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n341_), .B2(KEYINPUT20), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n319_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT20), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(new_n319_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT98), .B1(new_n350_), .B2(new_n334_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352_));
  AOI211_X1 g151(.A(new_n352_), .B(new_n335_), .C1(new_n346_), .C2(new_n349_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n336_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT91), .B1(new_n330_), .B2(new_n335_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n356_), .B(new_n334_), .C1(new_n321_), .C2(new_n329_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT92), .B1(new_n330_), .B2(new_n335_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT92), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n321_), .A2(new_n360_), .A3(new_n329_), .A4(new_n334_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n271_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n313_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n367_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT31), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n371_), .B(new_n376_), .Z(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n228_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n218_), .A3(new_n227_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT4), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n370_), .B1(new_n218_), .B2(new_n227_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n378_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n392_));
  OR3_X1    g191(.A1(new_n386_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n377_), .A2(new_n395_), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n270_), .A2(new_n354_), .A3(new_n364_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n330_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n341_), .A2(KEYINPUT20), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT96), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n316_), .A3(new_n343_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n348_), .B1(new_n404_), .B2(new_n319_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n401_), .B1(new_n405_), .B2(new_n398_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n398_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n350_), .A2(KEYINPUT97), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n400_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT33), .B(new_n390_), .C1(new_n386_), .C2(new_n392_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  INV_X1    g210(.A(new_n381_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(new_n383_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n380_), .A2(KEYINPUT94), .A3(new_n381_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n391_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n382_), .A2(new_n378_), .A3(new_n385_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n390_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n358_), .A2(new_n419_), .A3(new_n362_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n394_), .A2(KEYINPUT93), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT93), .B1(new_n394_), .B2(new_n421_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n270_), .B1(new_n409_), .B2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n268_), .A2(new_n269_), .A3(new_n395_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n354_), .A2(new_n427_), .A3(new_n364_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n397_), .B1(new_n429_), .B2(new_n377_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G229gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G1gat), .B(G8gat), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT76), .B(G15gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G22gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT76), .B(G15gat), .ZN(new_n438_));
  INV_X1    g237(.A(G22gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442_));
  INV_X1    g241(.A(G1gat), .ZN(new_n443_));
  INV_X1    g242(.A(G8gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT14), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n441_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n435_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n440_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n438_), .A2(new_n439_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n445_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT77), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n434_), .A3(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G29gat), .B(G36gat), .Z(new_n455_));
  XOR2_X1   g254(.A(G43gat), .B(G50gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n448_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n433_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n448_), .A2(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n457_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n457_), .B(KEYINPUT15), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n448_), .A3(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n432_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT82), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G169gat), .B(G197gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n475_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n471_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n478_));
  AOI211_X1 g277(.A(KEYINPUT81), .B(KEYINPUT82), .C1(new_n461_), .C2(new_n466_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G230gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT67), .B(G71gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G78gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G78gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n484_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n497_), .A2(new_n498_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  INV_X1    g304(.A(G92gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT9), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G85gat), .A3(G92gat), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n504_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n511_), .B(new_n504_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n503_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n507_), .A2(new_n508_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n500_), .A2(new_n502_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n519_), .B(new_n520_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  INV_X1    g326(.A(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n498_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n501_), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n521_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n520_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n518_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n517_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT66), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n517_), .B(new_n537_), .C1(new_n526_), .C2(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n494_), .A2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n532_), .A2(new_n533_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n519_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n532_), .A2(new_n518_), .A3(new_n533_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n494_), .A2(new_n539_), .B1(new_n541_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n490_), .A2(new_n493_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n536_), .A2(new_n550_), .A3(new_n538_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n551_), .A2(KEYINPUT70), .A3(new_n540_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT70), .B1(new_n551_), .B2(new_n540_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n483_), .B(new_n549_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n537_), .B1(new_n546_), .B2(new_n517_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n538_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n494_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n551_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  INV_X1    g358(.A(new_n483_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n551_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n550_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT68), .ZN(new_n565_));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  NAND4_X1  g369(.A1(new_n554_), .A2(new_n561_), .A3(new_n565_), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n559_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n574_));
  AOI211_X1 g373(.A(KEYINPUT68), .B(new_n483_), .C1(new_n557_), .C2(new_n551_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT72), .A3(new_n554_), .A4(new_n570_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n570_), .B1(new_n576_), .B2(new_n554_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n580_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(KEYINPUT73), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  AOI211_X1 g385(.A(new_n582_), .B(new_n579_), .C1(new_n573_), .C2(new_n577_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n580_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n482_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n458_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n548_), .A2(new_n464_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(KEYINPUT35), .B2(new_n594_), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n591_), .B(new_n595_), .C1(KEYINPUT35), .C2(new_n594_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n591_), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n597_), .B(new_n598_), .C1(new_n599_), .C2(new_n592_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n606_), .B(KEYINPUT36), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n596_), .B2(new_n600_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n609_), .A2(new_n612_), .A3(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n601_), .A2(new_n608_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n611_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G231gat), .ZN(new_n618_));
  INV_X1    g417(.A(G233gat), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n462_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n462_), .A2(new_n620_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n550_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n623_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n494_), .A3(new_n621_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT17), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n626_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT80), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n624_), .A2(new_n626_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT17), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n631_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT79), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(KEYINPUT79), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n637_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n617_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n431_), .A2(new_n590_), .A3(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT99), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(KEYINPUT99), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n443_), .A3(new_n395_), .A4(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n609_), .A2(new_n612_), .A3(KEYINPUT100), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT100), .B1(new_n609_), .B2(new_n612_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n431_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n590_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n646_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n395_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n651_), .A2(new_n652_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n653_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  NAND2_X1  g463(.A1(new_n354_), .A2(new_n364_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n649_), .A2(new_n444_), .A3(new_n665_), .A4(new_n650_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT101), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n444_), .B1(new_n659_), .B2(new_n665_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(KEYINPUT40), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n660_), .B2(new_n377_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n648_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n377_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n373_), .A3(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n679_), .A3(new_n682_), .ZN(G1326gat));
  XNOR2_X1  g482(.A(new_n270_), .B(KEYINPUT103), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n439_), .B1(new_n659_), .B2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT42), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n680_), .A2(new_n439_), .A3(new_n684_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1327gat));
  OR2_X1    g487(.A1(new_n613_), .A2(new_n616_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n430_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n681_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n617_), .B(new_n691_), .C1(new_n692_), .C2(new_n397_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n585_), .A2(new_n589_), .ZN(new_n695_));
  AND4_X1   g494(.A1(KEYINPUT104), .A2(new_n695_), .A3(new_n646_), .A4(new_n481_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n590_), .B2(new_n646_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n694_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n646_), .A3(new_n481_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n590_), .A2(KEYINPUT104), .A3(new_n646_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n701_), .A2(new_n702_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n704_));
  OAI21_X1  g503(.A(new_n698_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n661_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n658_), .A2(new_n430_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n646_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n656_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n661_), .A2(G29gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n706_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT106), .ZN(G1328gat));
  INV_X1    g513(.A(new_n665_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n710_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n698_), .B(new_n665_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n719_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT107), .B1(new_n719_), .B2(G36gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n718_), .B(KEYINPUT46), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n705_), .A2(new_n727_), .A3(new_n377_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n711_), .B2(new_n377_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1330gat));
  INV_X1    g532(.A(new_n270_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G50gat), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n705_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G50gat), .B1(new_n710_), .B2(new_n684_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1331gat));
  NOR3_X1   g538(.A1(new_n695_), .A2(new_n430_), .A3(new_n481_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n647_), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n395_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n695_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n646_), .A2(new_n481_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n746_), .A2(new_n657_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(new_n657_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n395_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n743_), .B1(new_n751_), .B2(new_n742_), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n715_), .A2(G64gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT110), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n741_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n665_), .A3(new_n749_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT111), .B(new_n755_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n681_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n741_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n750_), .A2(new_n681_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(G71gat), .ZN(new_n771_));
  AOI211_X1 g570(.A(KEYINPUT49), .B(new_n765_), .C1(new_n750_), .C2(new_n681_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  NAND3_X1  g572(.A1(new_n741_), .A2(new_n491_), .A3(new_n684_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n750_), .A2(new_n684_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G78gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT50), .B(new_n491_), .C1(new_n750_), .C2(new_n684_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1335gat));
  INV_X1    g578(.A(new_n694_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n695_), .A2(new_n708_), .A3(new_n481_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n661_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n740_), .A2(new_n709_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n505_), .A3(new_n395_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1336gat));
  OAI21_X1  g588(.A(G92gat), .B1(new_n784_), .B2(new_n715_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n506_), .A3(new_n665_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n497_), .A3(new_n681_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n681_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G99gat), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT113), .B(new_n528_), .C1(new_n783_), .C2(new_n681_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT114), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n798_), .B(new_n800_), .ZN(G1338gat));
  AOI21_X1  g600(.A(new_n498_), .B1(new_n783_), .B2(new_n734_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(KEYINPUT52), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n786_), .A2(G106gat), .A3(new_n270_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT115), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(new_n804_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n803_), .A2(new_n809_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n587_), .A2(new_n588_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n745_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n815_), .A3(new_n745_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n689_), .A3(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n814_), .A2(new_n689_), .A3(new_n816_), .A4(new_n818_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n549_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT55), .B1(new_n483_), .B2(KEYINPUT118), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT55), .B2(new_n483_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n570_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n830_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(KEYINPUT121), .A3(new_n832_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n467_), .A2(new_n477_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n463_), .A2(new_n839_), .A3(new_n465_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n433_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n459_), .A2(new_n460_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n433_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n838_), .B1(new_n844_), .B2(new_n477_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n578_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n824_), .B1(new_n836_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT58), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n824_), .B(new_n849_), .C1(new_n836_), .C2(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n617_), .A3(new_n850_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n476_), .A2(new_n480_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n833_), .A2(new_n835_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT119), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n853_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n581_), .A2(new_n845_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n656_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n859_), .B2(new_n656_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n851_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n646_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n823_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n665_), .A2(new_n734_), .A3(new_n661_), .A4(new_n377_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n867_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n863_), .A2(KEYINPUT123), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n851_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n646_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n873_), .B2(new_n823_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n481_), .B(new_n868_), .C1(new_n874_), .C2(new_n866_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G113gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n823_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n867_), .ZN(new_n878_));
  OR3_X1    g677(.A1(new_n878_), .A2(G113gat), .A3(new_n482_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1340gat));
  OAI211_X1 g679(.A(new_n744_), .B(new_n868_), .C1(new_n874_), .C2(new_n866_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G120gat), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n695_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n874_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(G1341gat));
  OAI211_X1 g685(.A(new_n708_), .B(new_n868_), .C1(new_n874_), .C2(new_n866_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G127gat), .ZN(new_n888_));
  OR3_X1    g687(.A1(new_n878_), .A2(G127gat), .A3(new_n646_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1342gat));
  OAI211_X1 g689(.A(new_n617_), .B(new_n868_), .C1(new_n874_), .C2(new_n866_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G134gat), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n878_), .A2(G134gat), .A3(new_n656_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1343gat));
  NOR4_X1   g693(.A1(new_n665_), .A2(new_n661_), .A3(new_n270_), .A4(new_n681_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n877_), .A2(new_n481_), .A3(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n877_), .A2(new_n744_), .A3(new_n895_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g698(.A1(new_n877_), .A2(new_n708_), .A3(new_n895_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(new_n656_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n877_), .A2(new_n212_), .A3(new_n903_), .A4(new_n895_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n877_), .A2(new_n617_), .A3(new_n895_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n212_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n665_), .A2(new_n396_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n684_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n823_), .B2(new_n864_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT22), .B(G169gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n481_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n859_), .A2(new_n656_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT57), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n859_), .A2(new_n656_), .A3(new_n860_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n708_), .B1(new_n917_), .B2(new_n851_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n481_), .B(new_n908_), .C1(new_n918_), .C2(new_n822_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n865_), .A2(KEYINPUT124), .A3(new_n481_), .A4(new_n908_), .ZN(new_n922_));
  AND4_X1   g721(.A1(new_n913_), .A2(new_n921_), .A3(G169gat), .A4(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n292_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n913_), .B1(new_n924_), .B2(new_n922_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n912_), .B1(new_n923_), .B2(new_n925_), .ZN(G1348gat));
  NOR3_X1   g725(.A1(new_n695_), .A2(new_n293_), .A3(new_n907_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n734_), .B(new_n928_), .C1(new_n873_), .C2(new_n823_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n910_), .B2(new_n744_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n932_), .A3(KEYINPUT125), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1349gat));
  INV_X1    g735(.A(new_n910_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n273_), .A2(new_n275_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n937_), .A2(new_n646_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n907_), .A2(new_n646_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n877_), .A2(new_n270_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n272_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n937_), .B2(new_n689_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n910_), .A2(new_n277_), .A3(new_n279_), .A4(new_n903_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1351gat));
  AND3_X1   g744(.A1(new_n665_), .A2(new_n427_), .A3(new_n377_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n877_), .A2(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947_), .B2(new_n481_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n877_), .A2(new_n946_), .ZN(new_n949_));
  INV_X1    g748(.A(G197gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n949_), .A2(new_n950_), .A3(new_n482_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n948_), .A2(new_n951_), .ZN(G1352gat));
  NOR2_X1   g751(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n744_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n954_), .B1(new_n947_), .B2(new_n957_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n949_), .A2(new_n956_), .A3(new_n953_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1353gat));
  AND2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  AOI211_X1 g761(.A(new_n961_), .B(new_n646_), .C1(KEYINPUT127), .C2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n877_), .A2(new_n946_), .A3(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n964_), .B(new_n965_), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n947_), .A2(new_n246_), .A3(new_n903_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G218gat), .B1(new_n949_), .B2(new_n689_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(G1355gat));
endmodule


