//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G85gat), .B(G92gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(KEYINPUT66), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT66), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .A4(new_n206_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n207_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT7), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT68), .A3(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n205_), .B1(new_n220_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n214_), .A2(new_n215_), .A3(new_n206_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n231_), .A2(KEYINPUT67), .B1(KEYINPUT7), .B2(new_n218_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n225_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n217_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n204_), .A2(KEYINPUT8), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n230_), .A2(KEYINPUT8), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT9), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n204_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G85gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT9), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n238_), .A2(new_n225_), .A3(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT10), .B(G99gat), .Z(new_n243_));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT10), .B(G99gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT64), .ZN(new_n247_));
  AOI21_X1  g046(.A(G106gat), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n246_), .B(new_n244_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n251_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n236_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT65), .B1(new_n251_), .B2(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n249_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n242_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT8), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n232_), .A2(new_n217_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n205_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n234_), .A2(new_n235_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT69), .B(new_n257_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G71gat), .B(G78gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT70), .Z(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n266_), .B2(KEYINPUT11), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(KEYINPUT70), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(KEYINPUT11), .A3(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n271_), .A2(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n254_), .A2(new_n276_), .A3(new_n262_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n254_), .A2(new_n276_), .A3(new_n262_), .A4(KEYINPUT71), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(KEYINPUT12), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n281_), .B1(new_n263_), .B2(new_n273_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n277_), .A2(KEYINPUT72), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n277_), .B2(new_n287_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n285_), .B(new_n286_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT73), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n277_), .A2(KEYINPUT72), .A3(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n283_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G120gat), .B(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(G204gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G176gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  AOI21_X1  g103(.A(new_n202_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n285_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n297_), .B1(new_n307_), .B2(new_n286_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n290_), .A2(KEYINPUT73), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n282_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n305_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n202_), .A3(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT13), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(KEYINPUT13), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT75), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT19), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT22), .B(G169gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n325_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT94), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G183gat), .ZN(new_n334_));
  INV_X1    g133(.A(G190gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n328_), .A2(new_n329_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT25), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G183gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(KEYINPUT25), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n331_), .B(KEYINPUT23), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n344_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT24), .B1(new_n324_), .B2(new_n325_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT93), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n346_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(KEYINPUT93), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n337_), .A2(new_n338_), .B1(new_n349_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G197gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(G204gat), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(KEYINPUT91), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT21), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n360_), .A2(KEYINPUT21), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n359_), .A2(new_n365_), .A3(KEYINPUT21), .A4(new_n360_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n356_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n340_), .B(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n341_), .A2(KEYINPUT82), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n341_), .A2(KEYINPUT82), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n343_), .A4(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n346_), .B(KEYINPUT84), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n333_), .B1(new_n374_), .B2(new_n347_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT85), .B1(new_n374_), .B2(new_n350_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377_));
  INV_X1    g176(.A(new_n350_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n353_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n345_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n328_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n367_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n323_), .B1(new_n368_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(new_n240_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT18), .B(G64gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n356_), .B2(new_n367_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n323_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n367_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n389_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT101), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n385_), .A2(new_n395_), .A3(KEYINPUT101), .A4(new_n389_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n368_), .A2(new_n384_), .A3(new_n323_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n327_), .A2(new_n325_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT94), .B1(new_n401_), .B2(new_n326_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n381_), .A3(new_n338_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n355_), .A2(new_n345_), .A3(new_n344_), .A4(new_n348_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n367_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT100), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT100), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(KEYINPUT20), .C1(new_n405_), .C2(new_n406_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n410_), .A3(new_n394_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n400_), .B1(new_n411_), .B2(new_n323_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n398_), .B(new_n399_), .C1(new_n412_), .C2(new_n389_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT27), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n407_), .A2(new_n323_), .A3(new_n393_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n390_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n392_), .B1(new_n416_), .B2(new_n383_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n389_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n389_), .B1(new_n385_), .B2(new_n395_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430_));
  INV_X1    g229(.A(G155gat), .ZN(new_n431_));
  INV_X1    g230(.A(G162gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n433_), .A2(new_n434_), .B1(KEYINPUT1), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n436_), .A2(new_n437_), .B1(KEYINPUT1), .B2(new_n435_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n436_), .A2(new_n437_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n428_), .B(new_n429_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT88), .B(KEYINPUT2), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n428_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT89), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n428_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n429_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT3), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n447_), .A2(new_n448_), .B1(new_n427_), .B2(KEYINPUT2), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n433_), .A2(new_n434_), .B1(G155gat), .B2(G162gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G228gat), .ZN(new_n455_));
  INV_X1    g254(.A(G233gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT92), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n440_), .B2(new_n452_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n454_), .B(new_n457_), .C1(new_n458_), .C2(new_n367_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n440_), .A2(new_n452_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n457_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n460_), .B(new_n453_), .C1(new_n406_), .C2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n424_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n424_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n464_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G22gat), .B(G50gat), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT92), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n467_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n380_), .A2(new_n382_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n481_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G127gat), .B(G134gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G113gat), .B(G120gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G227gat), .A2(G233gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT30), .B(G15gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT31), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n486_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n486_), .A2(new_n494_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n423_), .A2(new_n480_), .A3(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(new_n239_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n440_), .A2(new_n452_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n506_));
  INV_X1    g305(.A(new_n489_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n440_), .A2(new_n452_), .A3(new_n489_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT4), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n506_), .A3(new_n511_), .A4(new_n507_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n504_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n505_), .B(new_n489_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n504_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n503_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT96), .B(new_n489_), .C1(new_n440_), .C2(new_n452_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(KEYINPUT4), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n515_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n460_), .A2(new_n489_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n509_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n504_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n502_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n498_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n418_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n396_), .A3(KEYINPUT95), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n510_), .A2(new_n504_), .A3(new_n512_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n514_), .A2(new_n515_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n502_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT97), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(new_n503_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT98), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n502_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT97), .B1(KEYINPUT98), .B2(KEYINPUT33), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n535_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n526_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n385_), .A2(new_n395_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(KEYINPUT99), .Z(new_n549_));
  OAI22_X1  g348(.A1(new_n412_), .A2(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n480_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n479_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n476_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n423_), .A3(new_n546_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n497_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n527_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G43gat), .B(G50gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(G29gat), .B(G36gat), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT15), .Z(new_n570_));
  AOI22_X1  g369(.A1(new_n284_), .A2(new_n570_), .B1(new_n563_), .B2(new_n562_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n254_), .B2(new_n262_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n564_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n263_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n564_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n571_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT76), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n574_), .A2(new_n578_), .A3(new_n586_), .A4(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n581_), .B(KEYINPUT36), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n591_), .B2(KEYINPUT77), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n276_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G1gat), .B(G8gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT78), .ZN(new_n599_));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  INV_X1    g399(.A(G22gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G15gat), .A2(G22gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G1gat), .A2(G8gat), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n602_), .A2(new_n603_), .B1(KEYINPUT14), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n599_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n597_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT16), .B(G183gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n606_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n597_), .B(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(KEYINPUT17), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT79), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n559_), .A2(new_n595_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n570_), .A2(new_n614_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n606_), .A2(new_n575_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n606_), .B(new_n569_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n624_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT80), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n628_), .B2(new_n627_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT81), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n632_), .B(new_n633_), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n630_), .B(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n620_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n321_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n526_), .B(KEYINPUT102), .Z(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(G1gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OR3_X1    g440(.A1(new_n638_), .A2(KEYINPUT103), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT103), .B1(new_n638_), .B2(new_n641_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT38), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT95), .B1(new_n530_), .B2(new_n396_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n534_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT33), .B1(new_n537_), .B2(KEYINPUT98), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n531_), .B(new_n647_), .C1(new_n648_), .C2(new_n543_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n546_), .A2(new_n550_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n555_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n421_), .B1(new_n413_), .B2(KEYINPUT27), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n480_), .A2(new_n652_), .A3(new_n526_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n558_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n498_), .A2(new_n526_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n593_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n618_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n319_), .A3(new_n636_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT104), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G1gat), .B1(new_n662_), .B2(new_n546_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n644_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT38), .B1(new_n642_), .B2(new_n643_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1324gat));
  OAI21_X1  g465(.A(G8gat), .B1(new_n660_), .B2(new_n423_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n423_), .A2(G8gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n638_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n662_), .B2(new_n558_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n638_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n600_), .A3(new_n497_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(G1326gat));
  OR2_X1    g477(.A1(new_n555_), .A2(KEYINPUT106), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n555_), .A2(KEYINPUT106), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n601_), .B1(new_n661_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT42), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n676_), .A2(new_n601_), .A3(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT79), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n618_), .B(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(KEYINPUT111), .A3(new_n593_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n690_));
  INV_X1    g489(.A(new_n593_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n619_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n559_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n319_), .A3(new_n636_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n694_), .A2(G29gat), .A3(new_n546_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  INV_X1    g495(.A(new_n594_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n593_), .B(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n497_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n595_), .B(new_n702_), .C1(new_n703_), .C2(new_n527_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n705_));
  INV_X1    g504(.A(new_n700_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT108), .B(new_n706_), .C1(new_n559_), .C2(new_n698_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n656_), .A2(new_n708_), .A3(new_n702_), .A4(new_n595_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n701_), .A2(new_n705_), .A3(new_n707_), .A4(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n317_), .A2(new_n318_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n636_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n619_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n639_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n710_), .A2(new_n713_), .A3(KEYINPUT44), .A4(new_n619_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT110), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G29gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(KEYINPUT110), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n695_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n652_), .A3(new_n718_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n716_), .A2(KEYINPUT112), .A3(new_n652_), .A4(new_n718_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(G36gat), .A3(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n423_), .A2(G36gat), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n694_), .A2(KEYINPUT113), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT113), .B1(new_n694_), .B2(new_n729_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT45), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT114), .B(KEYINPUT46), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n728_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n558_), .A2(new_n483_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n716_), .A2(new_n718_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT115), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n716_), .A2(new_n743_), .A3(new_n718_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n483_), .B1(new_n694_), .B2(new_n558_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n749_), .A3(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1330gat));
  NAND3_X1  g550(.A1(new_n716_), .A2(new_n555_), .A3(new_n718_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G50gat), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n681_), .A2(G50gat), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT116), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n694_), .B2(new_n755_), .ZN(G1331gat));
  OR4_X1    g555(.A1(new_n321_), .A2(new_n636_), .A3(new_n619_), .A4(new_n657_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n526_), .A2(G57gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n319_), .A2(new_n636_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n620_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n639_), .ZN(new_n761_));
  OAI22_X1  g560(.A1(new_n757_), .A2(new_n758_), .B1(G57gat), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(G1332gat));
  OR3_X1    g562(.A1(new_n760_), .A2(G64gat), .A3(new_n423_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n757_), .A2(new_n423_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G64gat), .ZN(new_n767_));
  OAI211_X1 g566(.A(G64gat), .B(new_n765_), .C1(new_n757_), .C2(new_n423_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(G1333gat));
  OR3_X1    g569(.A1(new_n760_), .A2(G71gat), .A3(new_n558_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G71gat), .B1(new_n757_), .B2(new_n558_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT49), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(G71gat), .C1(new_n757_), .C2(new_n558_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n773_), .B2(new_n776_), .ZN(G1334gat));
  OR3_X1    g576(.A1(new_n760_), .A2(G78gat), .A3(new_n681_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G78gat), .B1(new_n757_), .B2(new_n681_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(G78gat), .C1(new_n757_), .C2(new_n681_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n780_), .B2(new_n783_), .ZN(G1335gat));
  AND2_X1   g583(.A1(new_n710_), .A2(new_n619_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n759_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(G85gat), .A3(new_n526_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n320_), .A2(new_n712_), .A3(new_n693_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n239_), .B1(new_n788_), .B2(new_n639_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n786_), .A2(G92gat), .A3(new_n652_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n240_), .B1(new_n788_), .B2(new_n423_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n793_), .B2(new_n792_), .ZN(G1337gat));
  OR2_X1    g594(.A1(new_n558_), .A2(new_n251_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT119), .B1(new_n788_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n786_), .A2(new_n497_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(G99gat), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n785_), .A2(new_n555_), .A3(new_n759_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(G106gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n802_), .B2(G106gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n555_), .A2(new_n213_), .ZN(new_n806_));
  OAI22_X1  g605(.A1(new_n804_), .A2(new_n805_), .B1(new_n788_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI221_X1 g608(.A(new_n809_), .B1(new_n788_), .B2(new_n806_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  NAND3_X1  g610(.A1(new_n698_), .A2(new_n712_), .A3(new_n688_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n319_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n319_), .B2(new_n813_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n624_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n634_), .B1(new_n626_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n819_), .A2(new_n820_), .B1(new_n623_), .B2(new_n818_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n630_), .A2(new_n635_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n313_), .A2(new_n314_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n299_), .A2(new_n304_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n636_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n291_), .B2(new_n298_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n285_), .B(new_n274_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n281_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n290_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n311_), .B1(new_n827_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT56), .B(new_n311_), .C1(new_n827_), .C2(new_n831_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n826_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n593_), .B1(new_n824_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n593_), .C1(new_n824_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n835_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n825_), .A3(new_n823_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n698_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n844_), .B2(new_n843_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n817_), .B1(new_n847_), .B2(new_n658_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n498_), .A3(new_n639_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n636_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  INV_X1    g650(.A(new_n848_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n498_), .A2(new_n639_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n851_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n688_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n817_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n854_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n636_), .B2(KEYINPUT122), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(KEYINPUT122), .B2(new_n861_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n850_), .B1(new_n860_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n319_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n849_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n854_), .A2(new_n859_), .A3(new_n321_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n849_), .B2(new_n688_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n618_), .A2(G127gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n860_), .B2(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n849_), .B2(new_n691_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n595_), .A2(G134gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT123), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n860_), .B2(new_n875_), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n848_), .A2(new_n497_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n639_), .A2(new_n480_), .A3(new_n652_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n712_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n425_), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n321_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n426_), .ZN(G1345gat));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n619_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT61), .B(G155gat), .Z(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  NOR3_X1   g685(.A1(new_n879_), .A2(new_n432_), .A3(new_n698_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n879_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n691_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n432_), .B2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n857_), .A2(new_n858_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n717_), .A2(new_n423_), .A3(new_n558_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n682_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895_), .B2(new_n712_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(KEYINPUT62), .B(G169gat), .C1(new_n895_), .C2(new_n712_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n895_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n636_), .A3(new_n327_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n899_), .A3(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n900_), .B2(new_n711_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n848_), .A2(new_n555_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n321_), .A2(new_n325_), .A3(new_n893_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n688_), .A3(new_n892_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n334_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n658_), .A2(new_n342_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT124), .B1(new_n895_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n895_), .A2(KEYINPUT124), .A3(new_n910_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1350gat));
  NAND4_X1  g713(.A1(new_n891_), .A2(new_n343_), .A3(new_n691_), .A4(new_n894_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n595_), .B(new_n894_), .C1(new_n856_), .C2(new_n817_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n916_), .A2(new_n917_), .A3(G190gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(G190gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n915_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT126), .B(new_n915_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n423_), .A2(new_n480_), .A3(new_n526_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n877_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n712_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n357_), .ZN(G1352gat));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n321_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n301_), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n877_), .A2(new_n618_), .A3(new_n925_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  XOR2_X1   g734(.A(KEYINPUT127), .B(G218gat), .Z(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n926_), .A2(new_n698_), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n926_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n691_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n940_), .B2(new_n937_), .ZN(G1355gat));
endmodule


