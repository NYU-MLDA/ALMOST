//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT81), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n205_), .B1(new_n209_), .B2(KEYINPUT82), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT82), .B2(new_n209_), .ZN(new_n211_));
  AND2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n208_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n204_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT4), .ZN(new_n229_));
  INV_X1    g028(.A(new_n227_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G1gat), .B(G29gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G85gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G57gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n235_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n234_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n240_), .B1(new_n245_), .B2(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT91), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT77), .B(G176gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT23), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n256_), .A2(KEYINPUT24), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT24), .A3(new_n248_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G190gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n252_), .A2(new_n255_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G211gat), .B(G218gat), .Z(new_n264_));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT86), .B1(G197gat), .B2(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n266_), .B(new_n267_), .C1(G204gat), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G204gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G197gat), .ZN(new_n273_));
  OAI221_X1 g072(.A(new_n273_), .B1(new_n272_), .B2(new_n270_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n265_), .A2(KEYINPUT86), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n264_), .A2(new_n275_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n263_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT76), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT25), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(KEYINPUT25), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n260_), .B(new_n281_), .C1(new_n282_), .C2(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n259_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n250_), .A2(new_n251_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n255_), .A2(new_n248_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT78), .ZN(new_n288_));
  INV_X1    g087(.A(new_n277_), .ZN(new_n289_));
  OAI211_X1 g088(.A(KEYINPUT20), .B(new_n278_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n289_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n263_), .B2(new_n277_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G8gat), .B(G36gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT95), .B1(new_n300_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  INV_X1    g107(.A(new_n306_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n308_), .B(new_n309_), .C1(new_n295_), .C2(new_n299_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n296_), .A2(new_n293_), .A3(new_n298_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n294_), .B2(new_n290_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n307_), .A2(new_n310_), .B1(new_n312_), .B2(new_n306_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n202_), .B1(new_n247_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n215_), .B2(new_n223_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n318_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n289_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI211_X1 g122(.A(new_n277_), .B(new_n323_), .C1(new_n317_), .C2(KEYINPUT84), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n317_), .A2(KEYINPUT84), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n321_), .A2(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G22gat), .B(G50gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n215_), .A2(new_n316_), .A3(new_n223_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n327_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT89), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT88), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n344_), .A3(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n326_), .A2(new_n346_), .A3(new_n337_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n340_), .A2(new_n343_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n326_), .B2(new_n337_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n326_), .A2(new_n337_), .A3(new_n346_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n247_), .A2(new_n313_), .A3(new_n202_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n315_), .A2(new_n348_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n246_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n312_), .A2(new_n305_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n312_), .A2(new_n305_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n228_), .A2(new_n235_), .A3(new_n231_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT94), .B1(new_n362_), .B2(new_n241_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT94), .A3(new_n241_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n365_));
  OAI221_X1 g164(.A(new_n361_), .B1(new_n355_), .B2(new_n246_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n354_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n312_), .A2(new_n305_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n371_), .B(KEYINPUT27), .C1(new_n305_), .C2(new_n300_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n247_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n352_), .A2(new_n348_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT79), .B(G15gat), .Z(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n288_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(new_n227_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  INV_X1    g182(.A(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n382_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n377_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n370_), .A2(new_n372_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n376_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n388_), .A2(new_n247_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n368_), .A2(new_n389_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT73), .B(G15gat), .ZN(new_n396_));
  INV_X1    g195(.A(G22gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G1gat), .ZN(new_n399_));
  INV_X1    g198(.A(G8gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT14), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G1gat), .B(G8gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G29gat), .B(G36gat), .Z(new_n406_));
  XOR2_X1   g205(.A(G43gat), .B(G50gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT74), .B1(new_n404_), .B2(new_n408_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G229gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT75), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n404_), .A2(new_n408_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(KEYINPUT75), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n413_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n415_), .A2(new_n421_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n395_), .A2(KEYINPUT97), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n376_), .A2(new_n394_), .A3(new_n390_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n352_), .A2(new_n348_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n247_), .A2(new_n313_), .A3(new_n202_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(new_n314_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n433_), .B(new_n435_), .C1(new_n358_), .C2(new_n366_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n388_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n431_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G230gat), .A2(G233gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT10), .B(G99gat), .Z(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G85gat), .A2(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(G99gat), .B2(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT6), .ZN(new_n458_));
  OAI221_X1 g257(.A(new_n454_), .B1(KEYINPUT9), .B2(new_n450_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n449_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(KEYINPUT6), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(G99gat), .A3(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n446_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n465_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n453_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n461_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT65), .B1(new_n456_), .B2(new_n458_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n469_), .A2(new_n470_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT66), .A3(new_n453_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n474_), .A2(KEYINPUT8), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n456_), .A2(new_n458_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n481_), .B(new_n453_), .C1(new_n482_), .C2(new_n471_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n460_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G71gat), .A2(G78gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(KEYINPUT11), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n488_), .B2(KEYINPUT11), .ZN(new_n491_));
  INV_X1    g290(.A(G64gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G57gat), .ZN(new_n493_));
  INV_X1    g292(.A(G57gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G64gat), .ZN(new_n495_));
  AND4_X1   g294(.A1(new_n490_), .A2(new_n493_), .A3(new_n495_), .A4(KEYINPUT11), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n495_), .A3(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT67), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n495_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n493_), .A2(new_n495_), .A3(new_n490_), .A4(KEYINPUT11), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n499_), .A2(new_n502_), .A3(new_n487_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n497_), .A2(new_n504_), .A3(KEYINPUT68), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n484_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT66), .B1(new_n478_), .B2(new_n453_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n483_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n460_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n509_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n444_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n484_), .B2(new_n509_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n444_), .B1(new_n484_), .B2(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n515_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n505_), .A2(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n517_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n530_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT13), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(KEYINPUT13), .A3(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT69), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT69), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n521_), .A2(new_n409_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n416_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n484_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT35), .B(new_n543_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n521_), .A2(new_n416_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n484_), .A2(new_n408_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT36), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n547_), .A2(new_n560_), .A3(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT37), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT37), .B1(new_n562_), .B2(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT72), .B1(new_n573_), .B2(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n404_), .B(new_n578_), .Z(new_n579_));
  AND2_X1   g378(.A1(new_n579_), .A2(new_n505_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n505_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  OR4_X1    g384(.A1(new_n577_), .A2(new_n580_), .A3(new_n581_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n509_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n579_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n579_), .A2(new_n587_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n585_), .B(KEYINPUT17), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n541_), .A2(new_n576_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n442_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT98), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n442_), .A2(new_n597_), .A3(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n374_), .A2(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n541_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n429_), .A3(new_n592_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606_));
  INV_X1    g405(.A(new_n561_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n557_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT100), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT100), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n395_), .A2(new_n606_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT101), .B1(new_n439_), .B2(new_n614_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n605_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n247_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G1gat), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n603_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n603_), .A2(KEYINPUT102), .A3(new_n620_), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1324gat));
  AOI211_X1 g425(.A(new_n373_), .B(new_n605_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT103), .B1(new_n627_), .B2(new_n400_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n618_), .A2(new_n390_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n631_), .A3(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  OAI211_X1 g432(.A(KEYINPUT103), .B(new_n633_), .C1(new_n627_), .C2(new_n400_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n596_), .A2(new_n598_), .A3(new_n400_), .A4(new_n390_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .A4(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  NAND2_X1  g440(.A1(new_n618_), .A2(new_n437_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n642_), .B2(G15gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n596_), .A2(new_n598_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n388_), .A2(G15gat), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n643_), .A2(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(G1326gat));
  NAND2_X1  g446(.A1(new_n618_), .A2(new_n376_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n648_), .A2(G22gat), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n648_), .B2(G22gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n376_), .A2(new_n397_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT106), .Z(new_n653_));
  OAI22_X1  g452(.A1(new_n650_), .A2(new_n651_), .B1(new_n645_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n615_), .A2(new_n592_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n442_), .A2(new_n604_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n247_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n541_), .A2(new_n440_), .A3(new_n592_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n395_), .B2(new_n576_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n439_), .A2(KEYINPUT43), .A3(new_n575_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665_));
  INV_X1    g464(.A(new_n658_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n395_), .A2(new_n659_), .A3(new_n576_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n575_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n669_), .B2(KEYINPUT44), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(KEYINPUT107), .A3(new_n663_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n664_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n247_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n657_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n672_), .B2(new_n390_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n373_), .A2(G36gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n656_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n442_), .A2(new_n604_), .A3(new_n655_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n680_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n682_), .A2(new_n678_), .A3(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n675_), .B1(new_n677_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n681_), .A2(new_n684_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n373_), .B(new_n664_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT46), .B(new_n687_), .C1(new_n688_), .C2(new_n676_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1329gat));
  NOR2_X1   g489(.A1(new_n388_), .A2(new_n384_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n672_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n656_), .A2(new_n437_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT109), .B(G43gat), .Z(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT47), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n672_), .A2(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n656_), .B2(new_n376_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n376_), .A2(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n672_), .B2(new_n702_), .ZN(G1331gat));
  NOR2_X1   g502(.A1(new_n439_), .A2(new_n429_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n576_), .A2(new_n593_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n541_), .A3(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT110), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n374_), .B1(new_n706_), .B2(KEYINPUT110), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n616_), .A2(new_n617_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n592_), .A2(new_n440_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n604_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(KEYINPUT111), .A3(new_n712_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n374_), .A2(new_n494_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n709_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n390_), .A3(new_n716_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G64gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G64gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n390_), .A2(new_n492_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n706_), .B2(new_n724_), .ZN(G1333gat));
  OR3_X1    g524(.A1(new_n706_), .A2(G71gat), .A3(new_n388_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n715_), .A2(new_n437_), .A3(new_n716_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G71gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1334gat));
  OR3_X1    g530(.A1(new_n706_), .A2(G78gat), .A3(new_n433_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n715_), .A2(new_n376_), .A3(new_n716_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(G78gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G78gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1335gat));
  NAND3_X1  g536(.A1(new_n541_), .A2(new_n440_), .A3(new_n593_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n374_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n541_), .A2(new_n655_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n704_), .A2(new_n742_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n743_), .A2(G85gat), .A3(new_n374_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n740_), .B2(new_n373_), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n743_), .A2(G92gat), .A3(new_n373_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1337gat));
  NOR2_X1   g547(.A1(new_n740_), .A2(new_n388_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n468_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n437_), .A2(new_n445_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n743_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1338gat));
  AOI21_X1  g554(.A(new_n446_), .B1(new_n739_), .B2(new_n376_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n376_), .A2(new_n446_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n758_), .A2(new_n759_), .B1(new_n743_), .B2(new_n760_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n418_), .A2(new_n420_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n413_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n766_), .B2(new_n765_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n412_), .A2(new_n414_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(new_n425_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n768_), .A2(new_n770_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n533_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n429_), .A2(new_n532_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n519_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n519_), .A2(new_n510_), .A3(new_n523_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n775_), .A2(KEYINPUT55), .B1(new_n444_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n524_), .A2(KEYINPUT114), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT114), .B1(new_n524_), .B2(new_n778_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n777_), .B(KEYINPUT115), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n529_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n774_), .B1(new_n787_), .B2(KEYINPUT116), .ZN(new_n788_));
  INV_X1    g587(.A(new_n785_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n522_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n516_), .A2(KEYINPUT12), .B1(new_n484_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n510_), .A2(new_n443_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n778_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n779_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT115), .B1(new_n796_), .B2(new_n777_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n529_), .B1(new_n789_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT56), .B(new_n529_), .C1(new_n789_), .C2(new_n797_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n773_), .B1(new_n788_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n764_), .B1(new_n804_), .B2(new_n614_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n801_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n787_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n798_), .A2(KEYINPUT116), .A3(new_n799_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n774_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n772_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n615_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n802_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n787_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n798_), .A2(KEYINPUT118), .A3(new_n799_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n771_), .A2(new_n532_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n800_), .A2(new_n814_), .A3(new_n802_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(KEYINPUT58), .A3(new_n817_), .A4(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n576_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n805_), .A2(new_n812_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n593_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n537_), .A2(new_n711_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n568_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n573_), .A2(KEYINPUT72), .A3(new_n569_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n575_), .A2(new_n832_), .A3(new_n826_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n831_), .A2(new_n833_), .B1(KEYINPUT113), .B2(KEYINPUT54), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n837_), .B(new_n834_), .C1(new_n824_), .C2(new_n593_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n392_), .A2(new_n374_), .A3(new_n388_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n429_), .ZN(new_n843_));
  AOI211_X1 g642(.A(KEYINPUT59), .B(new_n841_), .C1(new_n825_), .C2(new_n835_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n811_), .A2(new_n615_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n817_), .B(new_n818_), .C1(new_n815_), .C2(new_n787_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n575_), .B1(new_n846_), .B2(new_n813_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n845_), .A2(new_n764_), .B1(new_n847_), .B2(new_n822_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n592_), .B1(new_n848_), .B2(new_n812_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n837_), .B1(new_n849_), .B2(new_n834_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n825_), .A2(new_n835_), .A3(KEYINPUT119), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n840_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n844_), .B1(new_n853_), .B2(KEYINPUT59), .ZN(new_n854_));
  INV_X1    g653(.A(G113gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n429_), .B2(KEYINPUT120), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(KEYINPUT120), .B2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n843_), .B1(new_n854_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n604_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n842_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n604_), .B(new_n844_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n842_), .A2(new_n864_), .A3(new_n592_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n593_), .B(new_n844_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n842_), .A2(new_n868_), .A3(new_n614_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n575_), .B(new_n844_), .C1(new_n853_), .C2(KEYINPUT59), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1343gat));
  NAND3_X1  g670(.A1(new_n373_), .A2(new_n247_), .A3(new_n388_), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n433_), .B(new_n872_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n429_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n541_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n592_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT121), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT122), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n878_), .B(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(new_n883_), .A3(new_n614_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n873_), .A2(new_n576_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n883_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n825_), .A2(new_n835_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n376_), .A2(new_n394_), .A3(new_n373_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(new_n429_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G169gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n888_), .B(new_n889_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n891_), .ZN(new_n896_));
  OAI221_X1 g695(.A(new_n895_), .B1(KEYINPUT123), .B2(KEYINPUT62), .C1(new_n896_), .C2(new_n440_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n892_), .A2(new_n251_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n894_), .A2(new_n897_), .A3(KEYINPUT124), .A4(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1348gat));
  NOR2_X1   g702(.A1(new_n839_), .A2(new_n376_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n394_), .A2(new_n373_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n541_), .A2(G176gat), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n896_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n541_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n904_), .A2(new_n906_), .B1(new_n908_), .B2(new_n250_), .ZN(G1349gat));
  NOR3_X1   g708(.A1(new_n896_), .A2(new_n261_), .A3(new_n593_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(new_n592_), .A3(new_n905_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n280_), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n896_), .B2(new_n575_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n614_), .A2(new_n260_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n896_), .B2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT125), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n376_), .A2(new_n374_), .A3(new_n388_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n390_), .B1(new_n917_), .B2(KEYINPUT126), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(KEYINPUT126), .B2(new_n917_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT127), .B(new_n919_), .C1(new_n836_), .C2(new_n838_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924_), .B2(new_n429_), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n269_), .B(new_n440_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1352gat));
  AOI21_X1  g726(.A(KEYINPUT127), .B1(new_n852_), .B2(new_n919_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n923_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n541_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G204gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n924_), .A2(new_n272_), .A3(new_n541_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1353gat));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n592_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n924_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n937_), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n934_), .B(new_n939_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1354gat));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n924_), .A2(new_n942_), .A3(new_n614_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n575_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n942_), .B2(new_n944_), .ZN(G1355gat));
endmodule


