//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AOI22_X1  g005(.A1(KEYINPUT84), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(new_n204_), .ZN(new_n208_));
  OR3_X1    g007(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n202_), .B(new_n203_), .C1(new_n208_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT82), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n202_), .A2(new_n217_), .A3(KEYINPUT1), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n218_), .A4(new_n203_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G141gat), .B(G148gat), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT83), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n213_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G22gat), .B(G50gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n219_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n223_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n212_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n232_), .B2(KEYINPUT29), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT86), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n229_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G204gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT88), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(G204gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n242_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248_));
  AND2_X1   g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G211gat), .A2(G218gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT21), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n247_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n241_), .A2(G197gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n244_), .A2(G204gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n259_), .B(new_n260_), .C1(new_n258_), .C2(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n253_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n266_), .B(new_n264_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n268_), .A2(KEYINPUT90), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT90), .B1(new_n268_), .B2(new_n269_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n240_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT90), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G78gat), .B(G106gat), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n272_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n281_));
  OR2_X1    g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(G183gat), .B2(G190gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT23), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n285_), .B(KEYINPUT23), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n298_));
  OAI22_X1  g097(.A1(new_n295_), .A2(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OR3_X1    g098(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n288_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n294_), .A2(new_n299_), .A3(new_n300_), .A4(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n281_), .B1(new_n293_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G43gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n293_), .A2(new_n304_), .A3(new_n281_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(G43gat), .B1(new_n310_), .B2(new_n305_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G71gat), .B(G99gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT30), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G15gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  INV_X1    g121(.A(G120gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT79), .B(G113gat), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n325_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT31), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT78), .B1(new_n319_), .B2(new_n320_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n320_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n318_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n329_), .A2(KEYINPUT80), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(KEYINPUT80), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n332_), .A2(new_n335_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n339_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n331_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n225_), .A2(new_n328_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n324_), .B(new_n325_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n232_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT4), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n232_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT94), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n343_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n346_), .A2(KEYINPUT94), .A3(new_n348_), .A4(new_n350_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .A4(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n287_), .A2(new_n292_), .ZN(new_n368_));
  OR2_X1    g167(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(KEYINPUT91), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n373_));
  AOI21_X1  g172(.A(G176gat), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n304_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n253_), .A3(new_n262_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT20), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n293_), .A2(new_n304_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n253_), .B2(new_n262_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT92), .B(new_n367_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n264_), .B2(new_n378_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n367_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n375_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n263_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT18), .B(G64gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n384_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n377_), .A2(new_n367_), .A3(new_n379_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n386_), .A2(new_n389_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n367_), .B2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n365_), .B(new_n396_), .C1(new_n399_), .C2(new_n395_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n364_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n382_), .A2(new_n390_), .A3(new_n383_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n394_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n382_), .A2(new_n390_), .A3(new_n383_), .A4(new_n394_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n390_), .A4(new_n394_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n362_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n364_), .A2(new_n401_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n402_), .A2(new_n410_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n280_), .B(new_n342_), .C1(new_n400_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n417_), .A3(new_n409_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(KEYINPUT27), .C1(new_n394_), .C2(new_n399_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n418_), .A2(new_n277_), .A3(new_n279_), .A4(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT96), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n272_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n278_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n365_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n342_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n416_), .B1(new_n431_), .B2(KEYINPUT97), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n342_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n418_), .A2(new_n419_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n341_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n338_), .A2(new_n339_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n438_), .A2(new_n439_), .B1(new_n330_), .B2(new_n321_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n440_), .A3(new_n280_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n428_), .B1(new_n435_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n432_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(KEYINPUT12), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT6), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  OR3_X1    g248(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G85gat), .B(G92gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT8), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT9), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n452_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT64), .A3(G92gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n462_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n460_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT10), .B(G99gat), .Z(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n461_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n468_), .A2(new_n448_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n458_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n477_));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n446_), .B1(new_n474_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G230gat), .A2(G233gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n458_), .A2(new_n473_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n445_), .A2(KEYINPUT12), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n482_), .B(new_n483_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n483_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n474_), .A2(new_n481_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n484_), .A2(new_n485_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G204gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT5), .B(G176gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT68), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n494_), .B(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT74), .B(G1gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G8gat), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n513_), .B2(KEYINPUT14), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515_));
  AOI211_X1 g314(.A(KEYINPUT75), .B(new_n515_), .C1(new_n512_), .C2(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n510_), .B(new_n518_), .C1(new_n514_), .C2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT76), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n527_), .B(new_n528_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n529_));
  OAI22_X1  g328(.A1(new_n526_), .A2(new_n529_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n525_), .B(KEYINPUT15), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n520_), .A2(new_n521_), .A3(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n532_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n509_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n537_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n509_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n540_), .B(new_n541_), .C1(new_n537_), .C2(new_n536_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n506_), .A2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n444_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n522_), .B(new_n481_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G127gat), .B(G155gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT16), .B(G183gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT17), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n549_), .B1(new_n556_), .B2(new_n553_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n484_), .A2(new_n534_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n528_), .B2(new_n484_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT34), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(KEYINPUT35), .ZN(new_n564_));
  OR3_X1    g363(.A1(new_n560_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(KEYINPUT35), .A3(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(KEYINPUT72), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT69), .B(G190gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(KEYINPUT72), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT70), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n568_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n576_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT71), .B1(new_n567_), .B2(new_n574_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n584_), .B(KEYINPUT37), .C1(new_n585_), .C2(new_n580_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n558_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n546_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n512_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n365_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT38), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n576_), .A2(new_n580_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n558_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n546_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n428_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(G1324gat));
  OAI21_X1  g396(.A(G8gat), .B1(new_n595_), .B2(new_n437_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(KEYINPUT39), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(G8gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n588_), .A2(new_n603_), .A3(new_n436_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n599_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n602_), .A2(new_n606_), .A3(KEYINPUT40), .A4(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n595_), .B2(new_n440_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT41), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n588_), .A2(new_n315_), .A3(new_n342_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  XNOR2_X1  g414(.A(new_n280_), .B(KEYINPUT99), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G22gat), .B1(new_n595_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n588_), .A2(new_n621_), .A3(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n558_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n592_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n546_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n365_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n545_), .A2(new_n558_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n582_), .A2(new_n586_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n444_), .B2(new_n633_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT43), .B(new_n632_), .C1(new_n432_), .C2(new_n443_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(G29gat), .A3(new_n365_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n628_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n436_), .B(KEYINPUT102), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n627_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(new_n434_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n427_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n365_), .B1(new_n649_), .B2(new_n441_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n400_), .A2(new_n415_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n440_), .A3(new_n424_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n429_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n433_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n633_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n444_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n629_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n437_), .B1(new_n658_), .B2(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n638_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n647_), .B1(new_n660_), .B2(G36gat), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT101), .B(new_n643_), .C1(new_n659_), .C2(new_n638_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n646_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n646_), .B(KEYINPUT46), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1329gat));
  OAI21_X1  g466(.A(new_n307_), .B1(new_n626_), .B2(new_n440_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n638_), .A2(G43gat), .A3(new_n342_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n640_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g470(.A1(new_n641_), .A2(G50gat), .A3(new_n280_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n638_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n626_), .A2(new_n617_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n672_), .A2(new_n673_), .B1(G50gat), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT103), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n505_), .A2(new_n543_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n444_), .A2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(new_n558_), .A3(new_n633_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n365_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n678_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n594_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n365_), .A2(G57gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1332gat));
  INV_X1    g484(.A(new_n679_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n644_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n686_), .A2(G64gat), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G64gat), .B1(new_n682_), .B2(new_n687_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT48), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT48), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT104), .Z(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n682_), .B2(new_n440_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT49), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n440_), .A2(G71gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n686_), .B2(new_n696_), .ZN(G1334gat));
  OAI21_X1  g496(.A(G78gat), .B1(new_n682_), .B2(new_n617_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT50), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n617_), .A2(G78gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n686_), .B2(new_n700_), .ZN(G1335gat));
  NAND2_X1  g500(.A1(new_n681_), .A2(new_n625_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n365_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n677_), .A2(new_n558_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n428_), .A2(new_n462_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(new_n465_), .B1(new_n702_), .B2(new_n437_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT105), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n464_), .A2(new_n465_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n687_), .B1(new_n466_), .B2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n706_), .B2(new_n713_), .ZN(G1337gat));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n342_), .A2(new_n469_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n706_), .A2(new_n342_), .ZN(new_n717_));
  INV_X1    g516(.A(G99gat), .ZN(new_n718_));
  OAI221_X1 g517(.A(new_n715_), .B1(new_n702_), .B2(new_n716_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g519(.A(new_n705_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n280_), .B(new_n721_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT107), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n656_), .A2(new_n657_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n280_), .A4(new_n721_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(G106gat), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT52), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n723_), .A2(new_n729_), .A3(G106gat), .A4(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n703_), .A2(new_n470_), .A3(new_n280_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n735_), .A3(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(KEYINPUT54), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n506_), .A2(new_n543_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n587_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(KEYINPUT54), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT109), .Z(new_n743_));
  NOR2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n743_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n739_), .B(new_n745_), .C1(new_n587_), .C2(new_n740_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n494_), .A2(new_n498_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n489_), .A2(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT55), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n482_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n490_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n489_), .A2(KEYINPUT110), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n498_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n749_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n536_), .A2(KEYINPUT111), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n535_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n537_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n541_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n542_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(new_n542_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n502_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n759_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n592_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n772_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n757_), .A2(new_n758_), .A3(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(new_n748_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n756_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n498_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n779_), .B(new_n780_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n778_), .A2(new_n781_), .B1(new_n782_), .B2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(new_n768_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n765_), .A2(new_n766_), .A3(new_n542_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n748_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n756_), .A2(new_n498_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n782_), .A2(KEYINPUT58), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n786_), .A2(new_n792_), .A3(new_n793_), .A4(new_n780_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n633_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .A4(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n747_), .B1(new_n797_), .B2(new_n558_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n427_), .A2(new_n365_), .A3(new_n342_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n543_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT59), .B1(new_n799_), .B2(KEYINPUT116), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT57), .B1(new_n770_), .B2(new_n592_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n795_), .B2(new_n633_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n775_), .B1(new_n805_), .B2(KEYINPUT117), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n632_), .B1(new_n783_), .B2(new_n794_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n804_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n624_), .B1(new_n806_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n802_), .B(new_n803_), .C1(new_n810_), .C2(new_n747_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT118), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n796_), .A2(KEYINPUT117), .A3(new_n773_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n776_), .A3(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n558_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n747_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n800_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n543_), .A2(G113gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n801_), .B1(new_n823_), .B2(new_n824_), .ZN(G1340gat));
  OAI21_X1  g624(.A(new_n323_), .B1(new_n505_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT119), .B1(new_n323_), .B2(KEYINPUT60), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n800_), .B(new_n828_), .C1(new_n829_), .C2(new_n826_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n820_), .A2(new_n506_), .A3(new_n822_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n323_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n800_), .B2(new_n624_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n624_), .A2(G127gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n823_), .B2(new_n834_), .ZN(G1342gat));
  AOI21_X1  g634(.A(G134gat), .B1(new_n800_), .B2(new_n593_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n633_), .A2(G134gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n823_), .B2(new_n837_), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n440_), .A2(new_n280_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n798_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n365_), .A3(new_n687_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n544_), .ZN(new_n842_));
  INV_X1    g641(.A(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n505_), .ZN(new_n845_));
  INV_X1    g644(.A(G148gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n841_), .A2(new_n558_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(G162gat), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n841_), .A2(new_n851_), .A3(new_n632_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n841_), .B2(new_n592_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT120), .B(new_n851_), .C1(new_n841_), .C2(new_n592_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n687_), .A2(new_n365_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n342_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n617_), .B(new_n862_), .C1(new_n810_), .C2(new_n747_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n859_), .B(G169gat), .C1(new_n863_), .C2(new_n544_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n817_), .A2(new_n543_), .A3(new_n617_), .A4(new_n862_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n859_), .B1(new_n866_), .B2(G169gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n858_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n747_), .B1(new_n814_), .B2(new_n558_), .ZN(new_n869_));
  NOR4_X1   g668(.A1(new_n869_), .A2(new_n544_), .A3(new_n616_), .A4(new_n861_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n371_), .A2(new_n373_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n301_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(KEYINPUT62), .A3(new_n864_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n872_), .A3(new_n874_), .ZN(G1348gat));
  INV_X1    g674(.A(new_n863_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876_), .B2(new_n506_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n798_), .A2(new_n280_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n878_), .A2(G176gat), .A3(new_n506_), .A4(new_n862_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n880_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n877_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NOR2_X1   g682(.A1(new_n861_), .A2(new_n558_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G183gat), .B1(new_n878_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n863_), .A2(new_n558_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n296_), .A2(new_n295_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n863_), .B2(new_n632_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n593_), .B1(new_n298_), .B2(new_n297_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n863_), .B2(new_n890_), .ZN(G1351gat));
  NAND2_X1  g690(.A1(new_n840_), .A2(new_n860_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n244_), .B1(new_n892_), .B2(new_n544_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n840_), .A2(G197gat), .A3(new_n543_), .A4(new_n860_), .ZN(new_n896_));
  OAI211_X1 g695(.A(KEYINPUT123), .B(new_n244_), .C1(new_n892_), .C2(new_n544_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(G1352gat));
  NOR2_X1   g697(.A1(new_n892_), .A2(new_n505_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n241_), .ZN(G1353gat));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n558_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT124), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n892_), .B2(new_n903_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT126), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n904_), .B(new_n906_), .ZN(G1354gat));
  AND3_X1   g706(.A1(new_n840_), .A2(new_n593_), .A3(new_n860_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n633_), .A2(G218gat), .ZN(new_n909_));
  OAI22_X1  g708(.A1(new_n908_), .A2(G218gat), .B1(new_n892_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI221_X1 g711(.A(KEYINPUT127), .B1(new_n892_), .B2(new_n909_), .C1(new_n908_), .C2(G218gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


