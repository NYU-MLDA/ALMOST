//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT94), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(G204gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT92), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n207_), .A3(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G204gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(G197gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(new_n209_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT92), .B1(new_n215_), .B2(G197gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n218_), .B(new_n212_), .C1(new_n220_), .C2(new_n216_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT93), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n210_), .A2(new_n223_), .A3(new_n218_), .A4(new_n212_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n214_), .A2(KEYINPUT21), .B1(new_n225_), .B2(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT26), .ZN(new_n232_));
  INV_X1    g031(.A(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT25), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT98), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT23), .B1(new_n233_), .B2(new_n231_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G183gat), .A3(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n238_), .A2(KEYINPUT24), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n235_), .A2(KEYINPUT98), .A3(new_n240_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n237_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(KEYINPUT82), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(KEYINPUT23), .C1(new_n233_), .C2(new_n231_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n233_), .A2(new_n231_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n239_), .B(new_n252_), .C1(new_n257_), .C2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n250_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT20), .B1(new_n226_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n232_), .B1(new_n230_), .B2(KEYINPUT80), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(KEYINPUT25), .B2(new_n233_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n227_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n266_), .A2(new_n228_), .B1(new_n230_), .B2(KEYINPUT80), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n257_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n240_), .B(KEYINPUT81), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n248_), .A4(new_n270_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n236_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n272_));
  AOI21_X1  g071(.A(G176gat), .B1(new_n236_), .B2(KEYINPUT22), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT83), .B1(new_n236_), .B2(KEYINPUT22), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n247_), .A2(KEYINPUT84), .A3(new_n258_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT84), .B1(new_n247_), .B2(new_n258_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n239_), .B(new_n275_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n225_), .A2(new_n205_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n206_), .A2(KEYINPUT21), .A3(new_n213_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n204_), .B1(new_n262_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n204_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n226_), .A2(new_n261_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n284_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n289_), .B1(new_n284_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n202_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n262_), .A2(new_n283_), .A3(new_n204_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n292_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n284_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT27), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT104), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(KEYINPUT104), .A3(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n311_), .A2(KEYINPUT2), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n311_), .A2(KEYINPUT91), .A3(KEYINPUT2), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT91), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n309_), .B(new_n310_), .C1(new_n318_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n309_), .A2(new_n323_), .A3(KEYINPUT1), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n309_), .B2(KEYINPUT1), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n310_), .A4(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n319_), .B(KEYINPUT88), .Z(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n315_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n282_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT95), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G78gat), .B(G106gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n282_), .A2(new_n331_), .A3(new_n333_), .A4(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT28), .B1(new_n330_), .B2(KEYINPUT29), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n322_), .A2(new_n344_), .A3(new_n345_), .A4(new_n329_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT96), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT97), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT97), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n350_), .A2(KEYINPUT96), .A3(new_n354_), .A4(new_n351_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  INV_X1    g155(.A(new_n351_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n348_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n342_), .A2(new_n353_), .A3(new_n355_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n355_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n336_), .A2(new_n339_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n337_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G113gat), .B(G120gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n371_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(KEYINPUT87), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT31), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(KEYINPUT31), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n383_));
  OR3_X1    g182(.A1(new_n382_), .A2(G43gat), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(G43gat), .B1(new_n382_), .B2(new_n383_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n279_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT86), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n386_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n384_), .A2(new_n385_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n368_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n373_), .A2(new_n375_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n330_), .A2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n322_), .A2(new_n329_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT4), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n404_), .A2(KEYINPUT4), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT100), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n330_), .A2(new_n377_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n402_), .B2(new_n330_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(new_n409_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT101), .B(KEYINPUT0), .Z(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n308_), .A2(new_n400_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT105), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n297_), .A2(new_n303_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n426_), .A2(new_n422_), .A3(new_n368_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT32), .B(new_n289_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n284_), .A2(new_n294_), .A3(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n428_), .B(new_n430_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n295_), .A2(new_n296_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n418_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n409_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT102), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n412_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n435_), .B2(new_n412_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT103), .B1(new_n407_), .B2(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT103), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n439_), .B(new_n409_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n433_), .B(new_n437_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n419_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n410_), .A2(new_n413_), .A3(KEYINPUT33), .A4(new_n418_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n432_), .A2(new_n441_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n368_), .B1(new_n431_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n399_), .B1(new_n427_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT105), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n425_), .B1(new_n448_), .B2(new_n423_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT68), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n453_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n453_), .A2(new_n459_), .A3(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G71gat), .B(G78gat), .Z(new_n475_));
  NOR2_X1   g274(.A1(G57gat), .A2(G64gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G57gat), .A2(G64gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT69), .B1(new_n481_), .B2(new_n476_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n483_), .B2(KEYINPUT11), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n478_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n481_), .A2(new_n476_), .A3(KEYINPUT69), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT11), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT11), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n484_), .B1(new_n490_), .B2(new_n475_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT66), .B(G92gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT65), .B(G85gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n467_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n459_), .A2(new_n461_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT10), .B(G99gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n505_), .A2(KEYINPUT10), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(KEYINPUT10), .ZN(new_n507_));
  OAI211_X1 g306(.A(KEYINPUT64), .B(new_n504_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n500_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n498_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n499_), .B1(new_n498_), .B2(new_n509_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n474_), .B(new_n491_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT70), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n474_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n491_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(KEYINPUT12), .A3(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n522_), .A3(new_n513_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n515_), .A2(new_n520_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n513_), .B1(new_n518_), .B2(new_n512_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT5), .B(G176gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G120gat), .B(G148gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT72), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n524_), .A2(KEYINPUT72), .A3(new_n526_), .A4(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n512_), .A2(new_n522_), .A3(new_n513_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n522_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n516_), .A2(KEYINPUT12), .A3(new_n517_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT12), .B1(new_n516_), .B2(new_n517_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n525_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n530_), .B(KEYINPUT71), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n546_));
  AND2_X1   g345(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n535_), .B(new_n545_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n535_), .A2(new_n545_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n546_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G29gat), .B(G36gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT15), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560_));
  INV_X1    g359(.A(G1gat), .ZN(new_n561_));
  INV_X1    g360(.A(G8gat), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G1gat), .B(G8gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n557_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT77), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n566_), .B(new_n557_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n571_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT78), .B(G169gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G197gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n573_), .B(new_n581_), .C1(new_n572_), .C2(new_n576_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n550_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n449_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n516_), .A2(new_n559_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n516_), .A2(new_n557_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT35), .B(new_n590_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n590_), .A2(KEYINPUT35), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n516_), .B2(new_n559_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(KEYINPUT35), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n596_), .C1(new_n516_), .C2(new_n557_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT36), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n593_), .A2(new_n597_), .A3(new_n604_), .A4(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n588_), .B1(new_n606_), .B2(KEYINPUT74), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n566_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n517_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G211gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT16), .B(G183gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n610_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n610_), .A2(new_n615_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n603_), .A2(new_n620_), .A3(KEYINPUT37), .A4(new_n605_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n607_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT76), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n587_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n422_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n561_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n586_), .B(KEYINPUT106), .ZN(new_n628_));
  INV_X1    g427(.A(new_n399_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n445_), .A2(new_n431_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n368_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n426_), .A2(new_n368_), .A3(new_n422_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n423_), .B1(new_n634_), .B2(new_n424_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n423_), .A2(new_n424_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n606_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n619_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n628_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n641_), .B2(new_n422_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n627_), .A2(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(new_n308_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n624_), .A2(new_n562_), .A3(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n641_), .A2(new_n308_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(G8gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  NAND3_X1  g451(.A1(new_n624_), .A2(new_n387_), .A3(new_n629_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT107), .ZN(new_n654_));
  OAI21_X1  g453(.A(G15gat), .B1(new_n641_), .B2(new_n399_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1326gat));
  OAI21_X1  g456(.A(G22gat), .B1(new_n641_), .B2(new_n631_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n624_), .A2(new_n660_), .A3(new_n368_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n606_), .A2(new_n619_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n587_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G29gat), .B1(new_n664_), .B2(new_n625_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n607_), .A2(new_n621_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n637_), .B2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT43), .B(new_n667_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n639_), .B(new_n628_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n449_), .B2(new_n667_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n637_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n639_), .A4(new_n628_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n625_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n665_), .B1(new_n679_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n677_), .A3(new_n644_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n664_), .A2(new_n683_), .A3(new_n644_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT45), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n664_), .A2(new_n686_), .A3(new_n683_), .A4(new_n644_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(KEYINPUT46), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NAND2_X1  g492(.A1(new_n673_), .A2(new_n677_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n629_), .A2(G43gat), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n664_), .A2(new_n629_), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n694_), .A2(new_n695_), .B1(G43gat), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n664_), .B2(new_n368_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n368_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n678_), .B2(new_n700_), .ZN(G1331gat));
  NOR2_X1   g500(.A1(new_n449_), .A2(new_n585_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n550_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n640_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n422_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n702_), .B(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n703_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n625_), .A3(new_n623_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n705_), .ZN(G1332gat));
  OAI21_X1  g510(.A(G64gat), .B1(new_n704_), .B2(new_n308_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(new_n623_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n308_), .A2(G64gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n714_), .B2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n629_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n704_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(new_n629_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n721_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n714_), .A2(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n704_), .B2(new_n631_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT50), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n631_), .A2(G78gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n714_), .B2(new_n727_), .ZN(G1335gat));
  NOR3_X1   g527(.A1(new_n550_), .A2(new_n619_), .A3(new_n585_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n676_), .A2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(new_n422_), .A3(new_n494_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n708_), .A2(new_n703_), .A3(new_n663_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n464_), .B1(new_n732_), .B2(new_n422_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT110), .B(new_n464_), .C1(new_n732_), .C2(new_n422_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n731_), .B1(new_n735_), .B2(new_n736_), .ZN(G1336gat));
  NOR3_X1   g536(.A1(new_n730_), .A2(new_n308_), .A3(new_n493_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n709_), .A2(new_n644_), .A3(new_n663_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n465_), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n730_), .B2(new_n399_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n399_), .A2(new_n502_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n732_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n676_), .A2(new_n368_), .A3(new_n729_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n368_), .A2(new_n504_), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n747_), .A2(new_n748_), .B1(new_n732_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  OAI221_X1 g552(.A(new_n751_), .B1(new_n732_), .B2(new_n749_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(G113gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT72), .B1(new_n542_), .B2(new_n530_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n534_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n585_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n524_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n538_), .A2(KEYINPUT55), .A3(new_n541_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n520_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(G230gat), .A3(G233gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n544_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n544_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n759_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n575_), .A2(new_n570_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n582_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n584_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n535_), .B2(new_n545_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT57), .B(new_n606_), .C1(new_n770_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n544_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n544_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n585_), .B(new_n535_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n774_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n606_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n769_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n584_), .A2(new_n772_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT114), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n773_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n667_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n789_), .B(KEYINPUT114), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n785_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n785_), .A2(new_n788_), .A3(KEYINPUT58), .A4(new_n791_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n638_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT113), .B1(new_n801_), .B2(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n782_), .A2(new_n606_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n784_), .A2(new_n800_), .A3(new_n802_), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n639_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  INV_X1    g608(.A(new_n585_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n550_), .A2(new_n809_), .A3(new_n810_), .A4(new_n622_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT112), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n550_), .A2(new_n810_), .A3(new_n622_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n535_), .A2(new_n545_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n585_), .B1(new_n816_), .B2(new_n548_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n809_), .A4(new_n622_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n812_), .A2(new_n814_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n808_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n644_), .A2(new_n422_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n400_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n756_), .B1(new_n825_), .B2(new_n810_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n784_), .A2(new_n800_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n801_), .A2(KEYINPUT57), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n639_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n821_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n824_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n585_), .A2(G113gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT118), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n827_), .A2(new_n828_), .B1(new_n837_), .B2(new_n839_), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n836_), .B2(new_n550_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n825_), .B1(new_n842_), .B2(G120gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n550_), .A2(KEYINPUT60), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(G120gat), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(G1341gat));
  NOR2_X1   g645(.A1(new_n825_), .A2(new_n639_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(G127gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n836_), .A2(new_n639_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n825_), .B2(new_n606_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT120), .B(G134gat), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n829_), .A2(new_n668_), .A3(new_n835_), .A4(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT119), .B(new_n851_), .C1(new_n825_), .C2(new_n606_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n854_), .A2(new_n856_), .A3(new_n857_), .ZN(G1343gat));
  XNOR2_X1  g657(.A(KEYINPUT121), .B(G141gat), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n820_), .B1(new_n807_), .B2(new_n639_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n823_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n631_), .A2(new_n629_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n585_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n865_), .B2(new_n585_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n860_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n869_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n867_), .A3(new_n859_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n865_), .A2(new_n703_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g674(.A(new_n864_), .B1(new_n808_), .B2(new_n821_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n619_), .A3(new_n823_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n865_), .A2(new_n879_), .A3(new_n619_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1346gat));
  NAND3_X1  g683(.A1(new_n876_), .A2(new_n668_), .A3(new_n823_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G162gat), .ZN(new_n886_));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n865_), .A2(new_n887_), .A3(new_n638_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n308_), .A2(new_n625_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n399_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n368_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n833_), .A2(new_n585_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT125), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n833_), .A2(new_n900_), .A3(new_n585_), .A4(new_n897_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(G169gat), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n833_), .A2(new_n897_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n251_), .A3(new_n585_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n899_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n901_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NOR2_X1   g707(.A1(new_n896_), .A2(new_n237_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n822_), .A2(new_n631_), .A3(new_n703_), .A4(new_n909_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n833_), .A2(new_n703_), .A3(new_n897_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(G176gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT126), .ZN(G1349gat));
  AOI21_X1  g712(.A(new_n639_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n822_), .A2(new_n631_), .A3(new_n619_), .A4(new_n895_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n905_), .A2(new_n914_), .B1(new_n915_), .B2(new_n233_), .ZN(G1350gat));
  NAND4_X1  g715(.A1(new_n905_), .A2(new_n230_), .A3(new_n232_), .A4(new_n638_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n905_), .A2(new_n668_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n231_), .ZN(G1351gat));
  XNOR2_X1  g718(.A(new_n797_), .B(KEYINPUT115), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n920_), .A2(new_n794_), .B1(new_n777_), .B2(new_n783_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n806_), .A2(new_n802_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n619_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n863_), .B(new_n893_), .C1(new_n923_), .C2(new_n820_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n876_), .A2(new_n926_), .A3(new_n893_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928_), .B2(new_n585_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n876_), .B2(new_n893_), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n861_), .A2(KEYINPUT127), .A3(new_n864_), .A4(new_n894_), .ZN(new_n931_));
  OAI211_X1 g730(.A(G197gat), .B(new_n585_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n929_), .A2(new_n933_), .ZN(G1352gat));
  AOI21_X1  g733(.A(G204gat), .B1(new_n928_), .B2(new_n703_), .ZN(new_n935_));
  OAI211_X1 g734(.A(G204gat), .B(new_n703_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1353gat));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  OAI211_X1 g738(.A(new_n619_), .B(new_n939_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n639_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n941_));
  OR2_X1    g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(G1354gat));
  OAI211_X1 g743(.A(G218gat), .B(new_n668_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n606_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(G218gat), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(G1355gat));
endmodule


