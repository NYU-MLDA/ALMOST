//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT18), .B(G64gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206_));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT91), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n210_), .A4(KEYINPUT21), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G197gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G204gat), .ZN(new_n214_));
  INV_X1    g013(.A(G204gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(G197gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT21), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n207_), .B1(new_n217_), .B2(KEYINPUT89), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n219_), .A2(KEYINPUT89), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n206_), .B2(KEYINPUT21), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(KEYINPUT90), .A3(new_n220_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n221_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  AND3_X1   g026(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n234_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G183gat), .ZN(new_n242_));
  INV_X1    g041(.A(G183gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT25), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT26), .B(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n227_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n229_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT23), .A3(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .A4(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n234_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n240_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n226_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n230_), .A2(new_n255_), .A3(new_n232_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT82), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n242_), .A2(new_n244_), .A3(KEYINPUT79), .ZN(new_n266_));
  OR3_X1    g065(.A1(new_n243_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT26), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n257_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n230_), .A2(new_n273_), .A3(new_n255_), .A4(new_n232_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n265_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n239_), .A2(KEYINPUT83), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  AOI21_X1  g076(.A(G176gat), .B1(new_n235_), .B2(new_n236_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n234_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n252_), .A2(new_n231_), .A3(new_n249_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n226_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n259_), .A2(KEYINPUT20), .A3(new_n263_), .A4(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n275_), .A2(new_n281_), .A3(new_n212_), .A4(new_n225_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT20), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT95), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n226_), .A2(new_n258_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT95), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n285_), .A2(new_n289_), .A3(KEYINPUT20), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n262_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n291_), .B2(new_n262_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n205_), .B(new_n284_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT99), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT97), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n258_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT97), .B(new_n240_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(KEYINPUT20), .B(new_n283_), .C1(new_n300_), .C2(new_n226_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n262_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n287_), .A2(new_n263_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n205_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n296_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI211_X1 g106(.A(KEYINPUT99), .B(new_n205_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n295_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT27), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n284_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n305_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n295_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT87), .ZN(new_n318_));
  OR3_X1    g117(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  INV_X1    g119(.A(G141gat), .ZN(new_n321_));
  INV_X1    g120(.A(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n318_), .A2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n328_), .A2(KEYINPUT1), .B1(new_n321_), .B2(new_n322_), .ZN(new_n329_));
  OAI221_X1 g128(.A(new_n329_), .B1(new_n321_), .B2(new_n322_), .C1(KEYINPUT1), .C2(new_n317_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n327_), .A2(new_n334_), .A3(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  INV_X1    g140(.A(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  OR2_X1    g144(.A1(new_n336_), .A2(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n340_), .B(new_n345_), .C1(new_n348_), .C2(new_n339_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n345_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n340_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT98), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT98), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n355_), .B(new_n350_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n282_), .B(KEYINPUT30), .Z(new_n358_));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT84), .ZN(new_n362_));
  XOR2_X1   g161(.A(G15gat), .B(G43gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n358_), .A2(new_n359_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(new_n335_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n226_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(KEYINPUT92), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n375_), .A2(new_n226_), .B1(KEYINPUT92), .B2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n378_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n379_), .B(new_n382_), .C1(new_n378_), .C2(new_n380_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G22gat), .B(G50gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n387_), .B(new_n390_), .Z(new_n391_));
  OR3_X1    g190(.A1(new_n386_), .A2(KEYINPUT93), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n385_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n386_), .A2(new_n391_), .B1(KEYINPUT93), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n316_), .A2(new_n357_), .A3(new_n374_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n392_), .A2(new_n357_), .A3(new_n394_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n313_), .A2(new_n314_), .A3(new_n295_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n306_), .A2(new_n308_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n314_), .B1(new_n400_), .B2(new_n295_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT100), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n354_), .A2(new_n356_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n304_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n404_), .B(new_n406_), .C1(new_n405_), .C2(new_n312_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n350_), .B1(new_n348_), .B2(new_n339_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n339_), .B2(new_n338_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n313_), .A2(new_n295_), .A3(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n353_), .B(KEYINPUT33), .Z(new_n411_));
  OAI21_X1  g210(.A(new_n407_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n395_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT100), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n316_), .A2(new_n414_), .A3(new_n398_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n403_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n374_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n397_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G183gat), .B(G211gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G127gat), .B(G155gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT17), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(KEYINPUT17), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G57gat), .B(G64gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT11), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G71gat), .A2(G78gat), .ZN(new_n428_));
  OR2_X1    g227(.A1(G71gat), .A2(G78gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(new_n426_), .C2(KEYINPUT11), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT69), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(KEYINPUT69), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n427_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(G1gat), .ZN(new_n440_));
  INV_X1    g239(.A(G8gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G8gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n438_), .B(new_n445_), .Z(new_n446_));
  NAND2_X1  g245(.A1(G231gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  MUX2_X1   g247(.A(new_n424_), .B(new_n425_), .S(new_n448_), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT78), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n418_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT10), .B(G99gat), .Z(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT9), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n452_), .A2(new_n453_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n342_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT9), .A3(new_n455_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n457_), .A2(new_n458_), .A3(new_n461_), .A4(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n467_), .A2(KEYINPUT10), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(KEYINPUT10), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n453_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(new_n454_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(new_n465_), .A3(new_n461_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT65), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n467_), .A3(new_n453_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT66), .B1(new_n463_), .B2(new_n464_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n462_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(KEYINPUT67), .A3(new_n477_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n480_), .A2(new_n481_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n460_), .A2(KEYINPUT8), .A3(new_n455_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n462_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n455_), .B(new_n460_), .C1(new_n478_), .C2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n491_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n474_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G43gat), .B(G50gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(G29gat), .B(G36gat), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT15), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(KEYINPUT72), .A3(new_n504_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n503_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n490_), .A2(new_n466_), .A3(new_n473_), .A4(new_n495_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n488_), .A2(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n513_), .A2(KEYINPUT68), .A3(new_n466_), .A4(new_n473_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n507_), .A2(new_n508_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT35), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n507_), .A2(new_n508_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT34), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(KEYINPUT35), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G190gat), .B(G218gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT76), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n516_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n527_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n534_), .B(new_n533_), .C1(new_n527_), .C2(new_n536_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(KEYINPUT37), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT37), .B1(new_n539_), .B2(new_n540_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n451_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n512_), .A2(new_n514_), .A3(new_n438_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n498_), .A2(KEYINPUT12), .A3(new_n438_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n438_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n515_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT64), .Z(new_n554_));
  NAND4_X1  g353(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n547_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n438_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT5), .B(G176gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT71), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n560_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT13), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n445_), .B(new_n503_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n445_), .A2(new_n503_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n504_), .B2(new_n445_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  MUX2_X1   g373(.A(new_n571_), .B(new_n573_), .S(new_n574_), .Z(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n575_), .B(new_n578_), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n570_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n546_), .A2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n581_), .A2(G1gat), .A3(new_n357_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT38), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n539_), .A2(new_n540_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n418_), .A2(new_n450_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n580_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G1gat), .B1(new_n587_), .B2(new_n357_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(G1324gat));
  OAI21_X1  g388(.A(G8gat), .B1(new_n587_), .B2(new_n316_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT39), .ZN(new_n591_));
  INV_X1    g390(.A(new_n316_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n441_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n581_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(G1325gat));
  OAI21_X1  g395(.A(G15gat), .B1(new_n587_), .B2(new_n417_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT41), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n581_), .A2(G15gat), .A3(new_n417_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1326gat));
  OAI21_X1  g399(.A(G22gat), .B1(new_n587_), .B2(new_n395_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT42), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n395_), .A2(G22gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT102), .Z(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n581_), .B2(new_n604_), .ZN(G1327gat));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n606_), .B1(new_n418_), .B2(new_n544_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT43), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT43), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n606_), .B(new_n609_), .C1(new_n418_), .C2(new_n544_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n580_), .A2(new_n450_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(KEYINPUT44), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n618_), .A2(KEYINPUT104), .A3(new_n357_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT104), .B1(new_n618_), .B2(new_n357_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(G29gat), .A3(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n418_), .A2(new_n584_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n612_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n624_), .A2(G29gat), .A3(new_n357_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(G1328gat));
  NAND3_X1  g425(.A1(new_n616_), .A2(new_n592_), .A3(new_n617_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G36gat), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n624_), .A2(G36gat), .A3(new_n316_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1329gat));
  NAND2_X1  g436(.A1(new_n374_), .A2(G43gat), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n624_), .A2(new_n417_), .ZN(new_n639_));
  OAI22_X1  g438(.A1(new_n618_), .A2(new_n638_), .B1(G43gat), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g440(.A(G50gat), .B1(new_n618_), .B2(new_n395_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n395_), .A2(G50gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n624_), .B2(new_n643_), .ZN(G1331gat));
  INV_X1    g443(.A(new_n579_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n569_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n586_), .A2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT107), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT107), .ZN(new_n649_));
  AND4_X1   g448(.A1(G57gat), .A2(new_n648_), .A3(new_n404_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n646_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n545_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G57gat), .B1(new_n652_), .B2(new_n404_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1332gat));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n592_), .A3(new_n649_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G64gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT108), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT48), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n659_), .A3(G64gat), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n658_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n652_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n316_), .A2(G64gat), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT109), .Z(new_n665_));
  OAI22_X1  g464(.A1(new_n661_), .A2(new_n662_), .B1(new_n663_), .B2(new_n665_), .ZN(G1333gat));
  OR3_X1    g465(.A1(new_n663_), .A2(G71gat), .A3(new_n417_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n648_), .A2(new_n374_), .A3(new_n649_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT49), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G71gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G71gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1334gat));
  OR3_X1    g471(.A1(new_n663_), .A2(G78gat), .A3(new_n395_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n395_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n648_), .A2(new_n674_), .A3(new_n649_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT50), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(new_n676_), .A3(G78gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(G78gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(G1335gat));
  INV_X1    g478(.A(new_n450_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n651_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n611_), .A2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT110), .Z(new_n683_));
  OAI21_X1  g482(.A(G85gat), .B1(new_n683_), .B2(new_n357_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n622_), .A2(new_n680_), .A3(new_n651_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n342_), .A3(new_n404_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1336gat));
  OAI21_X1  g486(.A(G92gat), .B1(new_n683_), .B2(new_n316_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n685_), .A2(new_n459_), .A3(new_n592_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1337gat));
  OAI21_X1  g489(.A(G99gat), .B1(new_n682_), .B2(new_n417_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n685_), .A2(new_n452_), .A3(new_n374_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g493(.A1(new_n685_), .A2(new_n453_), .A3(new_n674_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n608_), .A2(new_n674_), .A3(new_n610_), .A4(new_n681_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT111), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n698_), .B2(G106gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n611_), .A2(KEYINPUT111), .A3(new_n674_), .A4(new_n681_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  AND4_X1   g501(.A1(new_n696_), .A2(new_n700_), .A3(G106gat), .A4(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n695_), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT53), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT53), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n695_), .C1(new_n699_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1339gat));
  INV_X1    g507(.A(KEYINPUT120), .ZN(new_n709_));
  INV_X1    g508(.A(G113gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n592_), .A2(new_n417_), .A3(new_n357_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT117), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n555_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n558_), .B1(new_n548_), .B2(new_n547_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(KEYINPUT55), .A3(new_n554_), .A4(new_n550_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n556_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n564_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n719_), .A2(new_n727_), .A3(KEYINPUT56), .A4(new_n564_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n720_), .A2(KEYINPUT114), .A3(new_n721_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n724_), .A2(new_n726_), .A3(new_n728_), .A4(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n573_), .A2(G229gat), .A3(G233gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n571_), .A2(new_n574_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n578_), .A3(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT112), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n555_), .A2(new_n559_), .A3(new_n565_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n730_), .A2(new_n731_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n731_), .B1(new_n730_), .B2(new_n739_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n740_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n712_), .B1(new_n744_), .B2(new_n544_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n730_), .A2(KEYINPUT58), .A3(new_n739_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n741_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n730_), .A2(new_n731_), .A3(new_n739_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n742_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n543_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n541_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(KEYINPUT117), .A3(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n745_), .A2(new_n746_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n722_), .A2(new_n725_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n645_), .A3(new_n737_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n568_), .B2(new_n736_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n584_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT118), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n761_), .A3(KEYINPUT57), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n680_), .B1(new_n753_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n544_), .A2(new_n579_), .A3(new_n569_), .A4(new_n680_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n395_), .B(new_n711_), .C1(new_n764_), .C2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n710_), .B1(new_n768_), .B2(new_n579_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(KEYINPUT59), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n579_), .A2(new_n710_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT119), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n709_), .B(new_n769_), .C1(new_n770_), .C2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n753_), .A2(new_n763_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n450_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n767_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT59), .A3(new_n395_), .A4(new_n711_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n768_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n772_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n769_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT120), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n783_), .ZN(G1340gat));
  AOI21_X1  g583(.A(new_n674_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n569_), .B2(G120gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n711_), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n768_), .A2(new_n779_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n768_), .A2(new_n779_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n570_), .B(new_n788_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G120gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n768_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n793_), .B2(new_n680_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n770_), .A2(new_n450_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g597(.A(G134gat), .B1(new_n793_), .B2(new_n585_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n770_), .A2(new_n544_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g600(.A1(new_n592_), .A2(new_n357_), .A3(new_n374_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n674_), .B(new_n802_), .C1(new_n764_), .C2(new_n767_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n579_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(new_n321_), .ZN(G1344gat));
  OR3_X1    g604(.A1(new_n803_), .A2(KEYINPUT122), .A3(new_n569_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT121), .B(G148gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT122), .B1(new_n803_), .B2(new_n569_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1345gat));
  NOR2_X1   g610(.A1(new_n803_), .A2(new_n450_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT123), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n812_), .B(new_n814_), .ZN(G1346gat));
  INV_X1    g614(.A(G162gat), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n803_), .A2(new_n816_), .A3(new_n544_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n803_), .A2(new_n584_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(new_n818_), .ZN(G1347gat));
  NOR3_X1   g618(.A1(new_n417_), .A2(new_n316_), .A3(new_n404_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n645_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n395_), .B(new_n821_), .C1(new_n764_), .C2(new_n767_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(KEYINPUT124), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT124), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(G169gat), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n785_), .A2(new_n237_), .A3(new_n821_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n823_), .A2(new_n824_), .A3(G169gat), .A4(new_n826_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n829_), .A3(new_n830_), .ZN(G1348gat));
  NAND2_X1  g630(.A1(new_n785_), .A2(new_n820_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n569_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(new_n238_), .ZN(G1349gat));
  NAND3_X1  g633(.A1(new_n785_), .A2(new_n680_), .A3(new_n820_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n245_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n243_), .B2(new_n835_), .ZN(G1350gat));
  OAI21_X1  g636(.A(G190gat), .B1(new_n832_), .B2(new_n544_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n585_), .A2(new_n246_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n832_), .B2(new_n839_), .ZN(G1351gat));
  NOR2_X1   g639(.A1(new_n316_), .A2(new_n374_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n398_), .B(new_n841_), .C1(new_n764_), .C2(new_n767_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n579_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n213_), .ZN(G1352gat));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n569_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n215_), .ZN(G1353gat));
  NOR2_X1   g645(.A1(new_n842_), .A2(new_n450_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n848_));
  OR2_X1    g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT63), .B(G211gat), .Z(new_n852_));
  AOI22_X1  g651(.A1(new_n850_), .A2(new_n851_), .B1(new_n847_), .B2(new_n852_), .ZN(G1354gat));
  OR3_X1    g652(.A1(new_n842_), .A2(G218gat), .A3(new_n584_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT127), .ZN(new_n855_));
  OAI21_X1  g654(.A(G218gat), .B1(new_n842_), .B2(new_n544_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1355gat));
endmodule


