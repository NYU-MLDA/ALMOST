//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n979_, new_n980_, new_n982_, new_n983_, new_n984_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n995_, new_n996_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G43gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(G43gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(G50gat), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n209_), .ZN(new_n211_));
  INV_X1    g010(.A(G50gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(new_n207_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G85gat), .B2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G85gat), .B2(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n222_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT65), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(KEYINPUT64), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT66), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n220_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT6), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT10), .B(G99gat), .Z(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n223_), .B1(new_n222_), .B2(new_n217_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n227_), .A2(KEYINPUT66), .A3(new_n228_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n219_), .A3(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n230_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT7), .ZN(new_n243_));
  INV_X1    g042(.A(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n237_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(new_n233_), .A3(new_n234_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n218_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT8), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n242_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n242_), .B2(new_n255_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n214_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT15), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n212_), .B1(new_n211_), .B2(new_n207_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n208_), .A2(G50gat), .A3(new_n209_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT15), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n242_), .A2(new_n255_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n205_), .B1(new_n259_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(KEYINPUT67), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n242_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n271_), .A2(new_n214_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(KEYINPUT71), .B2(new_n205_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n205_), .A2(KEYINPUT71), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(KEYINPUT72), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n259_), .A2(new_n267_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n268_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G134gat), .ZN(new_n282_));
  INV_X1    g081(.A(G162gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT36), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n276_), .A2(new_n279_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n268_), .ZN(new_n291_));
  AND4_X1   g090(.A1(KEYINPUT73), .A2(new_n288_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT73), .B1(new_n280_), .B2(new_n290_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n202_), .B(new_n287_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n280_), .A2(KEYINPUT73), .A3(new_n290_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(KEYINPUT75), .A3(new_n202_), .A4(new_n287_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n285_), .B(KEYINPUT74), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n280_), .B2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n296_), .A2(new_n302_), .B1(new_n304_), .B2(KEYINPUT37), .ZN(new_n305_));
  XOR2_X1   g104(.A(KEYINPUT76), .B(G22gat), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G15gat), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT76), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(G15gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319_));
  AND2_X1   g118(.A1(G57gat), .A2(G64gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G57gat), .A2(G64gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G57gat), .ZN(new_n323_));
  INV_X1    g122(.A(G64gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G57gat), .A2(G64gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT68), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n322_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G78gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G71gat), .ZN(new_n333_));
  INV_X1    g132(.A(G71gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G78gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n328_), .B(new_n336_), .C1(new_n322_), .C2(new_n327_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n318_), .B(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT77), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G155gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G183gat), .B(G211gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n347_), .A2(KEYINPUT17), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT79), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(KEYINPUT77), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n347_), .A2(KEYINPUT17), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n341_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT80), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n341_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n305_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT81), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(G183gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT25), .B(G183gat), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n362_), .B(new_n365_), .C1(new_n366_), .C2(new_n363_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n364_), .A2(KEYINPUT84), .A3(KEYINPUT85), .A4(G183gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT26), .B(G190gat), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT23), .ZN(new_n376_));
  OR2_X1    g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(KEYINPUT24), .A3(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n369_), .A2(KEYINPUT86), .A3(new_n371_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n379_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G71gat), .B(G99gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n383_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT87), .B(G15gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT30), .B(G43gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n400_), .A2(new_n404_), .A3(new_n402_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(G127gat), .A2(G134gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G127gat), .A2(G134gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(G113gat), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G127gat), .ZN(new_n413_));
  INV_X1    g212(.A(G134gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G113gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G127gat), .A2(G134gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n412_), .A2(new_n418_), .A3(G120gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(G120gat), .B1(new_n412_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n409_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .A4(new_n422_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(G197gat), .B(G204gat), .Z(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT21), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G155gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n283_), .A3(KEYINPUT89), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(G155gat), .B2(G162gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT90), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G155gat), .A3(G162gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n442_), .A3(KEYINPUT91), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447_));
  INV_X1    g246(.A(G141gat), .ZN(new_n448_));
  INV_X1    g247(.A(G148gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT3), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n445_), .A2(new_n446_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n442_), .A2(KEYINPUT1), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n439_), .A2(new_n441_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n437_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n448_), .A2(new_n449_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G141gat), .A2(G148gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n432_), .B1(new_n465_), .B2(KEYINPUT29), .ZN(new_n466_));
  INV_X1    g265(.A(G22gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n465_), .A2(KEYINPUT29), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT28), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n468_), .A2(new_n470_), .ZN(new_n473_));
  AND2_X1   g272(.A1(KEYINPUT92), .A2(G233gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(KEYINPUT92), .A2(G233gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(G228gat), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n212_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G78gat), .B(G106gat), .Z(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OR3_X1    g279(.A1(new_n472_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485_));
  INV_X1    g284(.A(new_n421_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n437_), .A2(new_n442_), .A3(KEYINPUT91), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT91), .B1(new_n437_), .B2(new_n442_), .ZN(new_n488_));
  AND4_X1   g287(.A1(new_n450_), .A2(new_n453_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n463_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n439_), .A2(new_n441_), .A3(new_n458_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n458_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n494_), .B2(new_n437_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT99), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n456_), .A2(new_n464_), .A3(new_n421_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n465_), .A2(KEYINPUT99), .A3(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n497_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n421_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n500_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT4), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT100), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n496_), .A2(KEYINPUT4), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n504_), .B1(new_n517_), .B2(new_n503_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G85gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n485_), .B1(new_n518_), .B2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G8gat), .B(G36gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G64gat), .B(G92gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n432_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G226gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT19), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n366_), .A2(KEYINPUT94), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n366_), .A2(KEYINPUT94), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n381_), .B1(new_n536_), .B2(new_n370_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n385_), .A2(KEYINPUT95), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n376_), .A2(new_n539_), .A3(new_n384_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n389_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n430_), .B(new_n431_), .Z(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT20), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n531_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n533_), .B(KEYINPUT93), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n383_), .A2(new_n432_), .A3(new_n390_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT98), .B(new_n530_), .C1(new_n545_), .C2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n530_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT98), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n546_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n537_), .A2(new_n541_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n548_), .B1(new_n558_), .B2(new_n432_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n533_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT86), .B1(new_n369_), .B2(new_n371_), .ZN(new_n561_));
  AOI211_X1 g360(.A(new_n373_), .B(new_n370_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n563_), .A2(new_n381_), .B1(new_n389_), .B2(new_n385_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n559_), .B(new_n560_), .C1(new_n564_), .C2(new_n432_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n530_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT97), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n557_), .A2(new_n565_), .A3(new_n569_), .A4(new_n566_), .ZN(new_n570_));
  AND4_X1   g369(.A1(new_n551_), .A2(new_n554_), .A3(new_n568_), .A4(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n515_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n502_), .A3(new_n514_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n501_), .A2(new_n503_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n524_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n516_), .B1(new_n513_), .B2(KEYINPUT100), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n510_), .B(new_n512_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n503_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n504_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT33), .A3(new_n523_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n525_), .A2(new_n571_), .A3(new_n575_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n566_), .A2(KEYINPUT32), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n557_), .A2(new_n583_), .A3(new_n565_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n533_), .B1(new_n531_), .B2(new_n544_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n547_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n583_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n578_), .A2(new_n579_), .A3(new_n524_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n524_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n584_), .B(new_n589_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n484_), .B1(new_n582_), .B2(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT27), .B(new_n567_), .C1(new_n587_), .C2(new_n566_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n554_), .A2(new_n568_), .A3(new_n551_), .A4(new_n570_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT27), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n591_), .A2(new_n592_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n484_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n427_), .B1(new_n594_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n426_), .A2(new_n600_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n605_), .A3(new_n483_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n599_), .B2(new_n483_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n338_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n266_), .A2(new_n611_), .A3(KEYINPUT12), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n271_), .B2(new_n340_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n269_), .A2(new_n270_), .A3(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n340_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n615_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n618_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT70), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT13), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT13), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n316_), .B(new_n214_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(G229gat), .A3(G233gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n316_), .A2(new_n214_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G229gat), .A2(G233gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n265_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n642_), .B(new_n643_), .C1(new_n644_), .C2(new_n316_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G169gat), .B(G197gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT82), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(G113gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(G141gat), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n645_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT83), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n639_), .A2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n361_), .A2(new_n610_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n600_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G1gat), .B1(new_n664_), .B2(new_n665_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n662_), .A2(new_n663_), .A3(new_n666_), .A4(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n280_), .A2(new_n286_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n602_), .B2(new_n609_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n639_), .A2(new_n655_), .A3(new_n359_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n663_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G1gat), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n361_), .A2(new_n663_), .A3(new_n610_), .A4(new_n661_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n667_), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n677_), .A2(new_n678_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n668_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n668_), .A2(new_n676_), .A3(new_n679_), .A4(KEYINPUT105), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1324gat));
  INV_X1    g483(.A(new_n599_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n671_), .A2(new_n685_), .A3(new_n672_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT106), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n671_), .A2(new_n688_), .A3(new_n685_), .A4(new_n672_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(G8gat), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT39), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(G8gat), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n662_), .A2(new_n309_), .A3(new_n685_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(KEYINPUT40), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1325gat));
  AND2_X1   g499(.A1(new_n671_), .A2(new_n672_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n426_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G15gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT107), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n705_), .A3(G15gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n662_), .A2(new_n312_), .A3(new_n426_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n704_), .A2(KEYINPUT41), .A3(new_n706_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n709_), .A2(new_n711_), .A3(new_n712_), .A4(new_n713_), .ZN(G1326gat));
  AOI21_X1  g513(.A(new_n467_), .B1(new_n701_), .B2(new_n484_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT42), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n662_), .A2(new_n467_), .A3(new_n484_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1327gat));
  NAND3_X1  g517(.A1(new_n638_), .A2(new_n654_), .A3(new_n359_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n597_), .A2(new_n598_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n483_), .A3(new_n595_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT102), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n603_), .B1(new_n722_), .B2(new_n606_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n599_), .A2(new_n484_), .A3(new_n600_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT33), .B1(new_n580_), .B2(new_n523_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n485_), .B(new_n524_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n573_), .A2(new_n524_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n597_), .B1(new_n574_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n502_), .B1(new_n572_), .B2(new_n514_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n523_), .B1(new_n730_), .B2(new_n504_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n588_), .B1(new_n731_), .B2(new_n590_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n727_), .A2(new_n729_), .B1(new_n732_), .B2(new_n584_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n724_), .B1(new_n733_), .B2(new_n484_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n723_), .B1(new_n734_), .B2(new_n427_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n296_), .A2(new_n302_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n304_), .A2(KEYINPUT37), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n735_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n610_), .A2(new_n740_), .A3(new_n305_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n719_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT44), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n663_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n742_), .A2(KEYINPUT44), .ZN(new_n745_));
  OAI21_X1  g544(.A(G29gat), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n610_), .A2(new_n670_), .A3(new_n359_), .A4(new_n661_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n600_), .A2(G29gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT109), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n747_), .B2(new_n749_), .ZN(G1328gat));
  INV_X1    g549(.A(G36gat), .ZN(new_n751_));
  INV_X1    g550(.A(new_n719_), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT43), .B(new_n738_), .C1(new_n602_), .C2(new_n609_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n740_), .B1(new_n610_), .B2(new_n305_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n599_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n751_), .B1(new_n757_), .B2(new_n743_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n670_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n602_), .B2(new_n609_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n599_), .A2(G36gat), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n359_), .A3(new_n661_), .A4(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT45), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT45), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n766_), .A2(new_n767_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n758_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n685_), .B1(new_n742_), .B2(KEYINPUT44), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n755_), .A2(new_n756_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G36gat), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n763_), .A2(new_n764_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n771_), .A2(new_n777_), .ZN(G1329gat));
  INV_X1    g577(.A(G43gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n747_), .B2(new_n427_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n743_), .A2(G43gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n426_), .B1(new_n742_), .B2(KEYINPUT44), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT47), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n782_), .B(new_n787_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1330gat));
  NAND2_X1  g588(.A1(new_n743_), .A2(new_n484_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G50gat), .B1(new_n790_), .B2(new_n745_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n484_), .A2(new_n212_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT112), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n747_), .B2(new_n793_), .ZN(G1331gat));
  AND4_X1   g593(.A1(new_n358_), .A2(new_n351_), .A3(new_n656_), .A4(new_n658_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n671_), .A2(new_n639_), .A3(new_n795_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n323_), .A3(new_n600_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n361_), .A2(new_n610_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n638_), .A2(new_n654_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n663_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n797_), .B1(new_n802_), .B2(new_n323_), .ZN(G1332gat));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n804_));
  INV_X1    g603(.A(new_n796_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n685_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(G64gat), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT48), .B(new_n324_), .C1(new_n805_), .C2(new_n685_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n685_), .A2(new_n324_), .ZN(new_n809_));
  OAI22_X1  g608(.A1(new_n807_), .A2(new_n808_), .B1(new_n800_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT113), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  OAI221_X1 g611(.A(new_n812_), .B1(new_n800_), .B2(new_n809_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1333gat));
  NAND3_X1  g613(.A1(new_n801_), .A2(new_n334_), .A3(new_n426_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G71gat), .B1(new_n796_), .B2(new_n427_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n816_), .A2(KEYINPUT49), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(KEYINPUT49), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n817_), .B2(new_n818_), .ZN(G1334gat));
  OAI21_X1  g618(.A(G78gat), .B1(new_n796_), .B2(new_n483_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT50), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n484_), .A2(new_n332_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n800_), .B2(new_n822_), .ZN(G1335gat));
  NAND3_X1  g622(.A1(new_n639_), .A2(new_n655_), .A3(new_n359_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n735_), .A2(new_n759_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G85gat), .B1(new_n825_), .B2(new_n663_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n824_), .B(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n600_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n826_), .B1(new_n830_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g630(.A(G92gat), .B1(new_n825_), .B2(new_n685_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n829_), .A2(new_n599_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g633(.A(G99gat), .B1(new_n829_), .B2(new_n427_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n825_), .A2(new_n236_), .A3(new_n426_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n825_), .A2(new_n237_), .A3(new_n484_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n828_), .B(new_n484_), .C1(new_n754_), .C2(new_n753_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n841_), .A3(G106gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n840_), .B2(G106gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT53), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n839_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1339gat));
  AOI21_X1  g647(.A(new_n614_), .B1(new_n613_), .B2(new_n617_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n618_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n613_), .A2(KEYINPUT55), .A3(new_n617_), .A4(new_n614_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT115), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n257_), .A2(new_n258_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT12), .B1(new_n854_), .B2(new_n611_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n266_), .A2(new_n611_), .A3(KEYINPUT12), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n619_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(KEYINPUT55), .A4(new_n614_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n851_), .A2(new_n853_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n627_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n654_), .A2(new_n628_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n640_), .A2(new_n643_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n643_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n642_), .B(new_n869_), .C1(new_n644_), .C2(new_n316_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n650_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n868_), .A2(KEYINPUT117), .A3(new_n650_), .A4(new_n870_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n653_), .A3(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n632_), .A2(new_n633_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n759_), .B1(new_n867_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880_));
  INV_X1    g679(.A(new_n875_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n852_), .B(new_n859_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n627_), .B1(new_n882_), .B2(new_n851_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n861_), .A2(new_n862_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n628_), .B1(new_n886_), .B2(KEYINPUT56), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n880_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n875_), .B1(new_n886_), .B2(KEYINPUT56), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n884_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(KEYINPUT58), .A4(new_n628_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n888_), .A2(new_n736_), .A3(new_n737_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n863_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n886_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n866_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n634_), .A2(new_n881_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(KEYINPUT57), .A3(new_n759_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n879_), .A2(new_n892_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n359_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n738_), .A2(new_n903_), .A3(new_n638_), .A4(new_n795_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n638_), .A2(new_n795_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT54), .B1(new_n905_), .B2(new_n305_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n600_), .B(new_n427_), .C1(new_n722_), .C2(new_n606_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(KEYINPUT118), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n901_), .A2(new_n359_), .B1(new_n906_), .B2(new_n904_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n909_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G113gat), .B1(new_n915_), .B2(new_n654_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n909_), .A2(KEYINPUT119), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT59), .B1(new_n909_), .B2(KEYINPUT119), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n908_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT59), .B1(new_n912_), .B2(new_n913_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n660_), .A2(new_n416_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n916_), .B1(new_n921_), .B2(new_n922_), .ZN(G1340gat));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n920_), .A3(new_n639_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n919_), .A2(new_n920_), .A3(KEYINPUT121), .A4(new_n639_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n926_), .A2(G120gat), .A3(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929_));
  AOI21_X1  g728(.A(G120gat), .B1(new_n639_), .B2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n910_), .B2(new_n914_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(G120gat), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n931_), .A2(KEYINPUT120), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT120), .B1(new_n931_), .B2(new_n932_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n928_), .B1(new_n933_), .B2(new_n934_), .ZN(G1341gat));
  INV_X1    g734(.A(new_n359_), .ZN(new_n936_));
  AOI21_X1  g735(.A(G127gat), .B1(new_n915_), .B2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n359_), .A2(new_n413_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n921_), .B2(new_n938_), .ZN(G1342gat));
  AOI21_X1  g738(.A(G134gat), .B1(new_n915_), .B2(new_n670_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n738_), .A2(new_n414_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n921_), .B2(new_n941_), .ZN(G1343gat));
  AOI21_X1  g741(.A(new_n426_), .B1(new_n902_), .B2(new_n907_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n663_), .A2(new_n484_), .A3(new_n599_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n654_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n639_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n936_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT61), .B(G155gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1346gat));
  AOI21_X1  g752(.A(G162gat), .B1(new_n946_), .B2(new_n670_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n944_), .A2(new_n283_), .A3(new_n945_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n305_), .B2(new_n955_), .ZN(G1347gat));
  NOR3_X1   g755(.A1(new_n603_), .A2(new_n484_), .A3(new_n599_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n908_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n654_), .A2(new_n387_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT122), .Z(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(KEYINPUT57), .B1(new_n899_), .B2(new_n759_), .ZN(new_n963_));
  AOI211_X1 g762(.A(new_n878_), .B(new_n670_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n936_), .B1(new_n965_), .B2(new_n892_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n904_), .A2(new_n906_), .ZN(new_n967_));
  OAI211_X1 g766(.A(new_n654_), .B(new_n957_), .C1(new_n966_), .C2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n969_));
  AND3_X1   g768(.A1(new_n968_), .A2(new_n969_), .A3(G169gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n968_), .B2(G169gat), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n962_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  OAI211_X1 g773(.A(KEYINPUT123), .B(new_n962_), .C1(new_n970_), .C2(new_n971_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(G1348gat));
  NOR2_X1   g775(.A1(new_n958_), .A2(new_n638_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(new_n388_), .ZN(G1349gat));
  NAND2_X1  g777(.A1(new_n959_), .A2(new_n936_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(G183gat), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n980_), .B1(new_n979_), .B2(new_n536_), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n958_), .B2(new_n738_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n670_), .A2(new_n371_), .ZN(new_n983_));
  XOR2_X1   g782(.A(new_n983_), .B(KEYINPUT124), .Z(new_n984_));
  OAI21_X1  g783(.A(new_n982_), .B1(new_n958_), .B2(new_n984_), .ZN(G1351gat));
  NOR3_X1   g784(.A1(new_n663_), .A2(new_n483_), .A3(new_n599_), .ZN(new_n986_));
  OAI211_X1 g785(.A(new_n427_), .B(new_n986_), .C1(new_n966_), .C2(new_n967_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n987_), .A2(KEYINPUT125), .ZN(new_n988_));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n943_), .A2(new_n989_), .A3(new_n986_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n655_), .B1(new_n988_), .B2(new_n990_), .ZN(new_n991_));
  XNOR2_X1  g790(.A(KEYINPUT126), .B(G197gat), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n991_), .B(new_n992_), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n988_), .A2(new_n990_), .ZN(new_n994_));
  AND3_X1   g793(.A1(new_n994_), .A2(G204gat), .A3(new_n639_), .ZN(new_n995_));
  AOI21_X1  g794(.A(G204gat), .B1(new_n994_), .B2(new_n639_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(new_n995_), .A2(new_n996_), .ZN(G1353gat));
  NAND2_X1  g796(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n989_), .B1(new_n943_), .B2(new_n986_), .ZN(new_n999_));
  INV_X1    g798(.A(new_n986_), .ZN(new_n1000_));
  NOR4_X1   g799(.A1(new_n912_), .A2(KEYINPUT125), .A3(new_n426_), .A4(new_n1000_), .ZN(new_n1001_));
  OAI211_X1 g800(.A(new_n936_), .B(new_n998_), .C1(new_n999_), .C2(new_n1001_), .ZN(new_n1002_));
  NOR2_X1   g801(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1003_));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004_));
  XNOR2_X1  g803(.A(new_n1003_), .B(new_n1004_), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1002_), .A2(new_n1005_), .ZN(new_n1006_));
  NAND2_X1  g805(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1007_));
  NAND4_X1  g806(.A1(new_n994_), .A2(new_n936_), .A3(new_n1007_), .A4(new_n998_), .ZN(new_n1008_));
  AND2_X1   g807(.A1(new_n1006_), .A2(new_n1008_), .ZN(G1354gat));
  AOI21_X1  g808(.A(G218gat), .B1(new_n994_), .B2(new_n670_), .ZN(new_n1010_));
  AOI21_X1  g809(.A(new_n738_), .B1(new_n988_), .B2(new_n990_), .ZN(new_n1011_));
  AOI21_X1  g810(.A(new_n1010_), .B1(G218gat), .B2(new_n1011_), .ZN(G1355gat));
endmodule


