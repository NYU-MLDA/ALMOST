//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT65), .ZN(new_n204_));
  INV_X1    g003(.A(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G57gat), .ZN(new_n206_));
  INV_X1    g005(.A(G57gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G64gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT65), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT11), .B1(new_n204_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G71gat), .B(G78gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n208_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n203_), .A2(KEYINPUT65), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n212_), .A3(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(KEYINPUT11), .B(new_n211_), .C1(new_n204_), .C2(new_n209_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G231gat), .A2(G233gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n221_), .A2(new_n222_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n223_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230_));
  INV_X1    g029(.A(G1gat), .ZN(new_n231_));
  INV_X1    g030(.A(G8gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT14), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G1gat), .B(G8gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n226_), .A2(new_n229_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n202_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n226_), .A2(new_n229_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(KEYINPUT67), .A3(new_n237_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G127gat), .B(G155gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT16), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G183gat), .B(G211gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n240_), .A2(new_n244_), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(KEYINPUT17), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT76), .B(new_n252_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT77), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n251_), .A2(new_n255_), .A3(new_n259_), .A4(new_n256_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G99gat), .A2(G106gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT6), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT9), .ZN(new_n268_));
  OR2_X1    g067(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(G85gat), .A2(G92gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(KEYINPUT9), .A3(new_n267_), .ZN(new_n274_));
  AND4_X1   g073(.A1(new_n266_), .A2(new_n268_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT7), .ZN(new_n277_));
  INV_X1    g076(.A(G99gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n270_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT64), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(new_n277_), .A3(new_n278_), .A4(new_n270_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n266_), .A2(new_n276_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n273_), .A2(new_n267_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT8), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n275_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(KEYINPUT8), .A3(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n221_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT66), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n283_), .A2(KEYINPUT8), .A3(new_n284_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT8), .B1(new_n283_), .B2(new_n284_), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n275_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n221_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n290_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n264_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT67), .B1(new_n219_), .B2(new_n220_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n219_), .A2(KEYINPUT67), .A3(new_n220_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n302_), .A2(new_n289_), .A3(KEYINPUT12), .A4(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n294_), .B2(new_n221_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n264_), .B1(new_n294_), .B2(new_n221_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G120gat), .B(G148gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G176gat), .B(G204gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n300_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n300_), .B2(new_n308_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n262_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT13), .A3(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT69), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n320_), .A3(KEYINPUT69), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G29gat), .B(G36gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G43gat), .B(G50gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n287_), .A2(new_n328_), .A3(new_n288_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT72), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G232gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(KEYINPUT35), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n328_), .B(KEYINPUT15), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n289_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(KEYINPUT35), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT71), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT73), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(KEYINPUT73), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n330_), .A2(KEYINPUT73), .A3(new_n339_), .A4(new_n336_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G190gat), .B(G218gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT74), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G134gat), .B(G162gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(KEYINPUT36), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n348_), .B(KEYINPUT36), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n342_), .A2(new_n343_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT37), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT37), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n335_), .A2(new_n242_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n236_), .B2(new_n328_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G229gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT78), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n236_), .B(new_n328_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(G229gat), .A3(G233gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G141gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G169gat), .B(G197gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n261_), .A2(new_n325_), .A3(new_n358_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375_));
  INV_X1    g174(.A(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G127gat), .ZN(new_n377_));
  INV_X1    g176(.A(G127gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G134gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G120gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G113gat), .ZN(new_n382_));
  INV_X1    g181(.A(G113gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G120gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n377_), .A2(new_n379_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n375_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT82), .B1(new_n380_), .B2(new_n385_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT83), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AND4_X1   g189(.A1(new_n377_), .A2(new_n379_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n377_), .A2(new_n379_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT82), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394_));
  INV_X1    g193(.A(new_n389_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n398_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n402_), .A2(KEYINPUT84), .A3(KEYINPUT85), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404_));
  INV_X1    g203(.A(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n399_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT80), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G71gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(new_n278_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT26), .B(G190gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(G176gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT24), .A3(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(KEYINPUT24), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n416_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G183gat), .ZN(new_n424_));
  INV_X1    g223(.A(G190gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT23), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G183gat), .A3(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(new_n417_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(KEYINPUT79), .A3(new_n428_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(KEYINPUT23), .C1(new_n424_), .C2(new_n425_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n424_), .A2(new_n425_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n430_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT81), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n441_), .B(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n413_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n402_), .A2(KEYINPUT84), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n413_), .A2(new_n445_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n409_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n408_), .B2(new_n403_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(KEYINPUT86), .A3(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT21), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT89), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT21), .ZN(new_n461_));
  AND2_X1   g260(.A1(G197gat), .A2(G204gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G197gat), .A2(G204gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n459_), .B(new_n461_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(G197gat), .A2(G204gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G197gat), .A2(G204gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT21), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G211gat), .B(G218gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT90), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n464_), .A2(new_n467_), .A3(new_n471_), .A4(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n462_), .A2(new_n463_), .A3(new_n458_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G211gat), .B(G218gat), .Z(new_n475_));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT91), .B1(new_n467_), .B2(new_n468_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT88), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(KEYINPUT1), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(KEYINPUT1), .B2(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  INV_X1    g288(.A(G141gat), .ZN(new_n490_));
  INV_X1    g289(.A(G148gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501_));
  XOR2_X1   g300(.A(G155gat), .B(G162gat), .Z(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n493_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n484_), .B1(new_n505_), .B2(KEYINPUT29), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n470_), .A2(new_n472_), .B1(new_n478_), .B2(new_n477_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT92), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n482_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n502_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT87), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n514_), .B2(new_n493_), .ZN(new_n515_));
  OAI211_X1 g314(.A(G228gat), .B(G233gat), .C1(new_n515_), .C2(new_n507_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G78gat), .B(G106gat), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT28), .B1(new_n505_), .B2(KEYINPUT29), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n514_), .A2(new_n521_), .A3(new_n522_), .A4(new_n493_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G22gat), .B(G50gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n520_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n518_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n509_), .A2(new_n516_), .A3(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n519_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n528_), .B1(new_n519_), .B2(new_n530_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n505_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n535_));
  OAI221_X1 g334(.A(new_n493_), .B1(new_n392_), .B2(new_n391_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(KEYINPUT97), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n505_), .A2(new_n390_), .A3(new_n396_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G225gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G1gat), .B(G29gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G85gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT0), .B(G57gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(KEYINPUT4), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n541_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n535_), .B2(KEYINPUT4), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n542_), .B(new_n546_), .C1(new_n548_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n540_), .A2(KEYINPUT4), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n535_), .A2(KEYINPUT4), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n549_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n546_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n537_), .A2(new_n556_), .A3(new_n539_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n549_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n534_), .A2(new_n551_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n429_), .A2(new_n561_), .A3(new_n438_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n429_), .A2(new_n438_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n432_), .B1(new_n563_), .B2(KEYINPUT94), .ZN(new_n564_));
  INV_X1    g363(.A(new_n437_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n562_), .A2(new_n564_), .B1(new_n423_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT20), .B1(new_n566_), .B2(new_n507_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n482_), .A2(new_n508_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n441_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G226gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT19), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT95), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  AOI221_X4 g373(.A(new_n481_), .B1(new_n477_), .B2(new_n478_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT92), .B1(new_n473_), .B2(new_n479_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n569_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT20), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n564_), .A2(new_n562_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n423_), .A2(new_n565_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n581_), .B2(new_n480_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n573_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G8gat), .B(G36gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT18), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G64gat), .B(G92gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n573_), .A2(KEYINPUT20), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n566_), .A2(new_n507_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n482_), .A2(new_n508_), .A3(new_n441_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n566_), .A2(KEYINPUT96), .A3(new_n507_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n574_), .A2(new_n585_), .A3(new_n589_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n589_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n599_));
  AOI211_X1 g398(.A(KEYINPUT95), .B(new_n573_), .C1(new_n577_), .C2(new_n582_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n550_), .B1(new_n540_), .B2(KEYINPUT4), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n549_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(KEYINPUT33), .A3(new_n546_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n560_), .A2(new_n597_), .A3(new_n601_), .A4(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n546_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n551_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n589_), .A2(KEYINPUT32), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n575_), .A2(new_n576_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n578_), .B1(new_n566_), .B2(new_n507_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n612_), .A2(new_n441_), .B1(new_n613_), .B2(KEYINPUT99), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(KEYINPUT99), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n573_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n577_), .A2(new_n573_), .A3(new_n582_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n574_), .A2(new_n585_), .A3(new_n596_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n609_), .B(new_n618_), .C1(new_n611_), .C2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n533_), .B1(new_n606_), .B2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n598_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n622_), .A2(new_n597_), .A3(KEYINPUT27), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT27), .B1(new_n601_), .B2(new_n597_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n551_), .B(new_n608_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n457_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n453_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n533_), .A2(new_n609_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n623_), .A2(new_n624_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n601_), .A2(new_n597_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT27), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n597_), .A3(KEYINPUT27), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT100), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n628_), .B(new_n629_), .C1(new_n631_), .C2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n374_), .B1(new_n627_), .B2(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(new_n231_), .A3(new_n609_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT101), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT101), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n643_), .A3(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n637_), .A2(new_n627_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n373_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n321_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n647_), .A2(new_n261_), .A3(new_n354_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n609_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n646_), .A3(new_n652_), .ZN(G1324gat));
  NOR2_X1   g452(.A1(new_n631_), .A2(new_n636_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n638_), .A2(new_n232_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G8gat), .B1(new_n650_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n650_), .B2(new_n457_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n457_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n638_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(new_n533_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G22gat), .B1(new_n650_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n638_), .A2(new_n673_), .A3(new_n533_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n258_), .A2(new_n260_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n649_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n358_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n647_), .B2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT43), .B(new_n358_), .C1(new_n637_), .C2(new_n627_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n677_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  AND4_X1   g484(.A1(G29gat), .A2(new_n684_), .A3(new_n609_), .A4(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n354_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n647_), .A2(new_n649_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n609_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n686_), .A2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n684_), .A2(new_n654_), .A3(new_n685_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n656_), .A2(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n691_), .A3(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT45), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(KEYINPUT46), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n684_), .A2(G43gat), .A3(new_n628_), .A4(new_n685_), .ZN(new_n706_));
  INV_X1    g505(.A(G43gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n692_), .B2(new_n457_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1330gat));
  AND4_X1   g510(.A1(G50gat), .A2(new_n684_), .A3(new_n533_), .A4(new_n685_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G50gat), .B1(new_n693_), .B2(new_n533_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1331gat));
  NAND3_X1  g513(.A1(new_n261_), .A2(new_n358_), .A3(new_n321_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT106), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n373_), .B1(new_n637_), .B2(new_n627_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(KEYINPUT106), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n717_), .A4(new_n718_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n609_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n207_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT108), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n726_), .A3(new_n207_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n325_), .A2(new_n676_), .A3(new_n687_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n717_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n717_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n651_), .A2(new_n207_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n725_), .A2(new_n727_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  NAND4_X1  g534(.A1(new_n720_), .A2(new_n722_), .A3(new_n205_), .A4(new_n654_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n654_), .A3(new_n732_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n736_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  NOR2_X1   g544(.A1(new_n457_), .A2(G71gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n720_), .A2(new_n722_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n733_), .A2(new_n667_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(G71gat), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G71gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n720_), .A2(new_n722_), .A3(new_n753_), .A4(new_n533_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n733_), .A2(new_n533_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G78gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT50), .B(new_n753_), .C1(new_n733_), .C2(new_n533_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  INV_X1    g558(.A(new_n325_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n690_), .A2(new_n717_), .A3(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(G85gat), .A3(new_n651_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n321_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n261_), .A2(new_n763_), .A3(new_n373_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT112), .B(new_n764_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n609_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n762_), .B1(new_n769_), .B2(G85gat), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT113), .B(new_n762_), .C1(new_n769_), .C2(G85gat), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1336gat));
  INV_X1    g573(.A(new_n761_), .ZN(new_n775_));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n654_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n767_), .A2(new_n654_), .A3(new_n768_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n776_), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n765_), .B2(new_n457_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n628_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n780_), .B(KEYINPUT114), .C1(new_n761_), .C2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n775_), .A2(new_n270_), .A3(new_n533_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n533_), .B(new_n764_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1339gat));
  NOR4_X1   g590(.A1(new_n654_), .A2(new_n533_), .A3(new_n651_), .A4(new_n453_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n373_), .A2(new_n315_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n294_), .A2(new_n305_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n219_), .A2(KEYINPUT67), .A3(new_n220_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n301_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n794_), .A2(new_n796_), .B1(new_n298_), .B2(new_n305_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT117), .A3(new_n291_), .A4(new_n296_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n304_), .A2(new_n306_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n297_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n263_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n797_), .A2(new_n803_), .A3(KEYINPUT55), .A4(new_n307_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .A4(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT118), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n308_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n313_), .B1(new_n802_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT56), .B(new_n313_), .C1(new_n802_), .C2(new_n809_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n793_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n360_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n360_), .A2(new_n815_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n362_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n364_), .A2(new_n362_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n370_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n372_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n319_), .B2(new_n315_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n354_), .B1(new_n814_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n354_), .C1(new_n814_), .C2(new_n822_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n812_), .A2(new_n813_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n821_), .A2(new_n316_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(KEYINPUT58), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n829_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n828_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n832_), .A2(new_n835_), .A3(new_n679_), .A4(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n261_), .B1(new_n827_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n321_), .A2(new_n373_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n261_), .A2(new_n358_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n261_), .A2(new_n358_), .A3(new_n842_), .A4(new_n839_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n792_), .B1(new_n838_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n383_), .A3(new_n373_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n847_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n848_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n837_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n676_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n847_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n792_), .C1(KEYINPUT122), .C2(KEYINPUT59), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n648_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n850_), .B1(new_n859_), .B2(new_n383_), .ZN(G1340gat));
  OAI21_X1  g659(.A(new_n381_), .B1(new_n763_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n849_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n381_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n325_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n381_), .ZN(G1341gat));
  NAND3_X1  g663(.A1(new_n849_), .A2(new_n378_), .A3(new_n261_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n676_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n378_), .ZN(G1342gat));
  NAND3_X1  g666(.A1(new_n849_), .A2(new_n376_), .A3(new_n687_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n358_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n376_), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n847_), .B1(new_n854_), .B2(new_n676_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n654_), .A2(new_n667_), .A3(new_n670_), .A4(new_n651_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n373_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n373_), .B(new_n872_), .C1(new_n838_), .C2(new_n847_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(G141gat), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n876_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n874_), .A2(new_n760_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n874_), .A2(new_n261_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  NAND2_X1  g686(.A1(new_n874_), .A2(new_n679_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G162gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n871_), .A2(G162gat), .A3(new_n354_), .A4(new_n873_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n890_), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n874_), .B2(new_n679_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT125), .B1(new_n895_), .B2(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n654_), .A2(new_n667_), .A3(new_n629_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n871_), .A2(new_n648_), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT22), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G169gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n417_), .B1(new_n900_), .B2(new_n898_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n871_), .A2(new_n899_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G176gat), .B1(new_n907_), .B2(new_n325_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n418_), .A3(new_n321_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n261_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n414_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n424_), .B2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n907_), .B2(new_n358_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n906_), .A2(new_n415_), .A3(new_n687_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n656_), .A2(new_n625_), .A3(new_n667_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n857_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n648_), .ZN(new_n919_));
  INV_X1    g718(.A(G197gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1352gat));
  NAND3_X1  g720(.A1(new_n857_), .A2(new_n760_), .A3(new_n917_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(G204gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(G204gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT127), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n925_), .B(new_n927_), .ZN(G1353gat));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AND2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n918_), .A2(new_n676_), .A3(new_n929_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n918_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n261_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(new_n929_), .ZN(G1354gat));
  OR3_X1    g733(.A1(new_n918_), .A2(G218gat), .A3(new_n354_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G218gat), .B1(new_n918_), .B2(new_n358_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


