//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n205_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n207_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G197gat), .A2(G204gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n210_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(new_n214_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT89), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT89), .B1(new_n229_), .B2(new_n234_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n222_), .B(new_n228_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n232_), .B(new_n233_), .C1(G183gat), .C2(G190gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n227_), .B(KEYINPUT90), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G169gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT91), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n239_), .B(new_n240_), .C1(new_n242_), .C2(G176gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n219_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n216_), .A2(new_n218_), .ZN(new_n245_));
  INV_X1    g044(.A(G183gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n246_), .B2(KEYINPUT78), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n220_), .B(new_n247_), .C1(new_n248_), .C2(KEYINPUT78), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n249_), .A2(new_n234_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(G169gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT22), .B1(new_n254_), .B2(KEYINPUT79), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(KEYINPUT22), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n255_), .C1(new_n256_), .C2(KEYINPUT79), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n227_), .A3(new_n239_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT20), .B1(new_n245_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n204_), .B1(new_n244_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n219_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(new_n245_), .B2(new_n259_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n261_), .B(new_n266_), .C1(new_n204_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT27), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT96), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n204_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n238_), .A2(new_n243_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n245_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n260_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n204_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n273_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(KEYINPUT96), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n265_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT99), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n244_), .A2(new_n204_), .A3(new_n260_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT96), .B1(new_n286_), .B2(new_n281_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n274_), .A2(new_n273_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT99), .A3(new_n265_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n272_), .B1(new_n285_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n278_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n267_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n265_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT27), .B1(new_n294_), .B2(new_n271_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n202_), .B1(new_n291_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n272_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT99), .B1(new_n289_), .B2(new_n265_), .ZN(new_n298_));
  AOI211_X1 g097(.A(new_n284_), .B(new_n266_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n295_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT100), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT82), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n305_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n259_), .B(KEYINPUT30), .Z(new_n310_));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G227gat), .A2(G233gat), .ZN(new_n312_));
  INV_X1    g111(.A(G71gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G15gat), .B(G43gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT80), .ZN(new_n317_));
  INV_X1    g116(.A(G99gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(G99gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n315_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(G99gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n318_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n314_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n311_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n310_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n323_), .A2(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n311_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n309_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n310_), .A2(new_n329_), .A3(new_n311_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n308_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT31), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n305_), .B(new_n306_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT84), .ZN(new_n348_));
  INV_X1    g147(.A(G141gat), .ZN(new_n349_));
  INV_X1    g148(.A(G148gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT2), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n351_), .A2(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(new_n356_), .A3(KEYINPUT85), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT85), .B1(new_n348_), .B2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n346_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n345_), .B1(KEYINPUT1), .B2(new_n343_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n349_), .A2(new_n350_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n363_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n308_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT92), .B(KEYINPUT4), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n346_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n348_), .A2(new_n356_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n374_), .B2(new_n357_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n339_), .B1(new_n375_), .B2(new_n365_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n308_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(KEYINPUT4), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT93), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  INV_X1    g190(.A(new_n378_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n380_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n382_), .B(new_n388_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n391_), .B(new_n388_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT98), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT98), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n391_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n388_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n399_), .B1(new_n402_), .B2(new_n396_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n342_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n375_), .A2(new_n365_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n360_), .A2(new_n366_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n411_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n406_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT28), .B1(new_n411_), .B2(KEYINPUT29), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n405_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(KEYINPUT87), .A3(new_n416_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n245_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(G78gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G106gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n421_), .B(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n420_), .A2(new_n427_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n303_), .A2(new_n404_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n394_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT33), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n294_), .A2(new_n271_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n376_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n389_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n380_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n438_), .B2(new_n378_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n394_), .A2(new_n432_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n434_), .A2(new_n440_), .A3(KEYINPUT95), .A4(new_n442_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n266_), .A2(KEYINPUT32), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n292_), .A2(new_n293_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n289_), .B2(new_n447_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n395_), .A2(new_n397_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n430_), .B1(new_n403_), .B2(new_n398_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n291_), .A2(new_n295_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n451_), .A2(new_n430_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n342_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n431_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G15gat), .B(G22gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT76), .B(G1gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(G8gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G8gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n457_), .B(new_n462_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G29gat), .B(G36gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT15), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n472_), .A2(new_n464_), .A3(new_n465_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n466_), .B(new_n471_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(new_n478_), .B2(new_n476_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n477_), .B(new_n482_), .C1(new_n478_), .C2(new_n476_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT77), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n456_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G231gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n466_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n313_), .A2(KEYINPUT67), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT67), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G71gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n494_), .A3(new_n423_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G57gat), .B(G64gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(KEYINPUT11), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT67), .B(G71gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n423_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT68), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G64gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G57gat), .ZN(new_n502_));
  INV_X1    g301(.A(G57gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n493_), .A2(G71gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n313_), .A2(KEYINPUT67), .ZN(new_n509_));
  OAI21_X1  g308(.A(G78gat), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n503_), .A2(G64gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n501_), .A2(G57gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n510_), .A2(new_n513_), .A3(new_n514_), .A4(new_n495_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n500_), .A2(new_n507_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n507_), .B1(new_n500_), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n491_), .B(new_n518_), .Z(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT16), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n524_), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n519_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT64), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT64), .ZN(new_n535_));
  OR2_X1    g334(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n425_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(G85gat), .B(G92gat), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n538_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(G85gat), .ZN(new_n551_));
  INV_X1    g350(.A(G92gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n545_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n540_), .A2(KEYINPUT66), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT6), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n558_), .A3(new_n539_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT7), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n318_), .A3(new_n425_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n539_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n555_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n553_), .A2(new_n545_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n562_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n543_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n554_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n550_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n469_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n550_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n571_), .B(new_n573_), .C1(KEYINPUT35), .C2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT74), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(KEYINPUT36), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n586_));
  INV_X1    g385(.A(new_n578_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n576_), .B(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n588_), .B2(KEYINPUT75), .ZN(new_n589_));
  AND4_X1   g388(.A1(KEYINPUT75), .A2(new_n579_), .A3(new_n580_), .A4(new_n586_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT37), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n585_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n530_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n507_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n506_), .A2(new_n505_), .B1(new_n498_), .B2(new_n423_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n514_), .B1(new_n597_), .B2(new_n510_), .ZN(new_n598_));
  AND4_X1   g397(.A1(new_n514_), .A2(new_n510_), .A3(new_n513_), .A4(new_n495_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n500_), .A2(new_n507_), .A3(new_n515_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n572_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT70), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n570_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT70), .B1(new_n607_), .B2(new_n604_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n601_), .A3(new_n572_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n609_), .A2(KEYINPUT69), .A3(KEYINPUT12), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT12), .B1(new_n609_), .B2(KEYINPUT69), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n606_), .A2(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n604_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G120gat), .B(G148gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT72), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n609_), .A2(KEYINPUT69), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT12), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n609_), .A2(KEYINPUT69), .A3(KEYINPUT12), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n603_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n607_), .A2(KEYINPUT70), .A3(new_n604_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n613_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT72), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n620_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n622_), .A2(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n625_), .A2(new_n626_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n619_), .B1(new_n635_), .B2(new_n613_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n595_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n489_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n403_), .A2(new_n398_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n458_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n486_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT101), .ZN(new_n649_));
  INV_X1    g448(.A(new_n591_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n456_), .A2(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n649_), .A2(new_n529_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n644_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n645_), .A2(new_n646_), .B1(new_n654_), .B2(G1gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n646_), .B2(new_n645_), .ZN(G1324gat));
  INV_X1    g455(.A(G8gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n303_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n652_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT39), .Z(new_n660_));
  INV_X1    g459(.A(new_n643_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n652_), .B2(new_n455_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n661_), .A2(new_n669_), .A3(new_n455_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n430_), .B(KEYINPUT103), .Z(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n652_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n674_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT104), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n643_), .B2(new_n679_), .ZN(G1327gat));
  OR2_X1    g479(.A1(new_n649_), .A2(new_n530_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n592_), .A2(new_n594_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n451_), .A2(new_n430_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n452_), .A2(new_n453_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n455_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n303_), .A2(new_n404_), .A3(new_n430_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n682_), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n682_), .B1(new_n456_), .B2(new_n683_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n681_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n681_), .B2(new_n691_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n693_), .A2(G29gat), .A3(new_n653_), .A4(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n530_), .A2(new_n650_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n647_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n489_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n644_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(G29gat), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT105), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n693_), .A2(new_n658_), .A3(new_n694_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G36gat), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n698_), .A2(G36gat), .A3(new_n303_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT45), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n693_), .A2(G43gat), .A3(new_n455_), .A4(new_n694_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n698_), .A2(new_n342_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g513(.A(new_n698_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G50gat), .B1(new_n715_), .B2(new_n675_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n693_), .A2(new_n694_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n430_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n717_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n486_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n456_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n647_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n595_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n653_), .ZN(new_n727_));
  OR4_X1    g526(.A1(new_n488_), .A2(new_n651_), .A3(new_n647_), .A4(new_n529_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n644_), .A2(KEYINPUT106), .ZN(new_n730_));
  MUX2_X1   g529(.A(KEYINPUT106), .B(new_n730_), .S(G57gat), .Z(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n729_), .B2(new_n731_), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n728_), .B2(new_n303_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n501_), .A3(new_n658_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n728_), .B2(new_n342_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n313_), .A3(new_n455_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  AOI21_X1  g539(.A(new_n423_), .B1(new_n729_), .B2(new_n675_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT50), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n726_), .A2(new_n423_), .A3(new_n675_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1335gat));
  NAND3_X1  g543(.A1(new_n722_), .A2(new_n723_), .A3(new_n696_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n551_), .A3(new_n653_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT43), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(KEYINPUT107), .A3(new_n688_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n530_), .A2(new_n486_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n723_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT108), .B1(new_n753_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n755_), .C1(new_n749_), .C2(new_n752_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n757_), .A2(new_n759_), .A3(new_n644_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n747_), .B1(new_n760_), .B2(new_n551_), .ZN(G1336gat));
  OAI21_X1  g560(.A(new_n552_), .B1(new_n745_), .B2(new_n303_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT109), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n757_), .A2(new_n759_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n303_), .A2(new_n552_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1337gat));
  OAI211_X1 g565(.A(new_n746_), .B(new_n455_), .C1(new_n534_), .C2(new_n537_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT110), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n757_), .A2(new_n759_), .A3(new_n342_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n318_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n768_), .C1(new_n769_), .C2(new_n318_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  NAND2_X1  g573(.A1(new_n751_), .A2(new_n688_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n755_), .A2(new_n430_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n425_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n746_), .A2(new_n425_), .A3(new_n718_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n642_), .B2(new_n487_), .ZN(new_n785_));
  AND4_X1   g584(.A1(new_n784_), .A2(new_n647_), .A3(new_n487_), .A4(new_n724_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  INV_X1    g588(.A(new_n476_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n470_), .A2(new_n475_), .A3(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n483_), .B(new_n791_), .C1(new_n478_), .C2(new_n790_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n485_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT111), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n485_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n632_), .B1(new_n631_), .B2(new_n620_), .ZN(new_n798_));
  NOR4_X1   g597(.A1(new_n635_), .A2(KEYINPUT72), .A3(new_n613_), .A4(new_n619_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n602_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n635_), .A2(KEYINPUT55), .B1(new_n801_), .B2(new_n604_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n612_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n619_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n635_), .A2(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n612_), .A2(new_n803_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n605_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n619_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n800_), .B1(new_n807_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n789_), .B(new_n683_), .C1(new_n814_), .C2(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n485_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n795_), .B1(new_n485_), .B2(new_n792_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n622_), .B2(new_n633_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n612_), .A2(new_n803_), .B1(new_n810_), .B2(new_n605_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n806_), .B(new_n620_), .C1(new_n822_), .C2(new_n808_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n619_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n789_), .B1(new_n827_), .B2(new_n683_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n817_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n486_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n807_), .B2(new_n813_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n820_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n834_), .B2(new_n591_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n650_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n529_), .B1(new_n829_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n788_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n658_), .A2(new_n718_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n644_), .A2(new_n342_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n487_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT114), .B1(new_n817_), .B2(new_n828_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n807_), .A2(new_n813_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT58), .B1(new_n851_), .B2(new_n821_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n683_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT113), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n816_), .A4(new_n815_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n836_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n835_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n857_), .B(new_n830_), .C1(new_n834_), .C2(new_n591_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n850_), .A2(new_n856_), .A3(new_n859_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n529_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n842_), .B1(new_n862_), .B2(new_n788_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n849_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n787_), .B1(new_n861_), .B2(new_n529_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT116), .B(KEYINPUT59), .C1(new_n866_), .C2(new_n842_), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n845_), .B(new_n848_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n866_), .A2(new_n721_), .A3(new_n842_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT115), .B1(new_n869_), .B2(G113gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n788_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n842_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n486_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n846_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n783_), .B1(new_n868_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n865_), .A2(new_n867_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n844_), .A3(new_n847_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n870_), .A2(new_n875_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(KEYINPUT117), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n647_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n863_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n845_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n886_), .A2(new_n723_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n883_), .ZN(G1341gat));
  AOI21_X1  g687(.A(G127gat), .B1(new_n863_), .B2(new_n530_), .ZN(new_n889_));
  INV_X1    g688(.A(G127gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n530_), .B2(KEYINPUT118), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(KEYINPUT118), .B2(new_n890_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n886_), .B2(new_n892_), .ZN(G1342gat));
  AOI21_X1  g692(.A(G134gat), .B1(new_n863_), .B2(new_n591_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n683_), .A2(G134gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT119), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n886_), .B2(new_n896_), .ZN(G1343gat));
  NAND4_X1  g696(.A1(new_n303_), .A2(new_n653_), .A3(new_n718_), .A4(new_n342_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT120), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n871_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n721_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n349_), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n647_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n350_), .ZN(G1345gat));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n529_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  INV_X1    g706(.A(G162gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n900_), .B2(new_n650_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT121), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n900_), .A2(new_n908_), .A3(new_n853_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1347gat));
  AOI21_X1  g711(.A(new_n675_), .B1(new_n788_), .B2(new_n838_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n303_), .A2(new_n653_), .A3(new_n342_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n486_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n916_), .A3(G169gat), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n915_), .A2(new_n242_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n915_), .B2(G169gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n913_), .A2(new_n723_), .A3(new_n914_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n866_), .A2(new_n718_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n723_), .A2(new_n914_), .A3(G176gat), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n253_), .A2(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  AND2_X1   g724(.A1(new_n914_), .A2(new_n530_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G183gat), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n221_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n913_), .B2(new_n929_), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n913_), .A2(new_n683_), .A3(new_n914_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT122), .B1(new_n931_), .B2(G190gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n913_), .A2(new_n914_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n591_), .A2(new_n220_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT123), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n933_), .A2(new_n934_), .B1(new_n935_), .B2(new_n937_), .ZN(G1351gat));
  NAND3_X1  g737(.A1(new_n658_), .A2(new_n452_), .A3(new_n342_), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n866_), .A2(new_n207_), .A3(new_n721_), .A4(new_n939_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n940_), .A2(KEYINPUT124), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(KEYINPUT124), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n866_), .A2(new_n939_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943_), .B2(new_n486_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n941_), .A2(new_n942_), .A3(new_n944_), .ZN(G1352gat));
  NOR3_X1   g744(.A1(new_n866_), .A2(new_n647_), .A3(new_n939_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n206_), .A2(new_n208_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(G204gat), .B2(new_n946_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT125), .ZN(G1353gat));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951_));
  INV_X1    g750(.A(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n530_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT126), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n943_), .A2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n951_), .A2(new_n952_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n955_), .B(new_n956_), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n943_), .B2(new_n591_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n683_), .A2(G218gat), .ZN(new_n959_));
  XOR2_X1   g758(.A(new_n959_), .B(KEYINPUT127), .Z(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n943_), .B2(new_n960_), .ZN(G1355gat));
endmodule


