//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT25), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G190gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT77), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n213_), .A2(new_n214_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n205_), .B2(new_n209_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n217_), .A2(new_n219_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(new_n215_), .B2(new_n216_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n206_), .A2(new_n208_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT76), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n222_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n235_), .B(new_n237_), .C1(new_n226_), .C2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n204_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G71gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n241_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT31), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT79), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n249_), .B2(new_n248_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G99gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n252_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT80), .B1(new_n256_), .B2(KEYINPUT1), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(G155gat), .A4(G162gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(KEYINPUT1), .ZN(new_n261_));
  OR2_X1    g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n257_), .A2(new_n260_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G141gat), .B(G148gat), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  INV_X1    g065(.A(G141gat), .ZN(new_n267_));
  INV_X1    g066(.A(G148gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n269_), .A2(new_n272_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n262_), .A2(new_n256_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n265_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT29), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G228gat), .A2(G233gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT83), .Z(new_n281_));
  NOR2_X1   g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n283_));
  INV_X1    g082(.A(G197gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(G204gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G204gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(new_n293_), .A3(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(G197gat), .B2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n289_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n286_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(G204gat), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n282_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT21), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n292_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n279_), .A2(new_n281_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(KEYINPUT85), .ZN(new_n305_));
  INV_X1    g104(.A(new_n279_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n304_), .B1(new_n307_), .B2(new_n281_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G78gat), .B(G106gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n309_), .B(new_n304_), .C1(new_n307_), .C2(new_n281_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n313_));
  OR3_X1    g112(.A1(new_n278_), .A2(KEYINPUT29), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n278_), .B2(KEYINPUT29), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G22gat), .B(G50gat), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n317_), .A3(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT82), .B1(new_n319_), .B2(new_n320_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n311_), .B(new_n312_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n308_), .A2(KEYINPUT86), .A3(new_n309_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n309_), .A2(KEYINPUT86), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n304_), .C1(new_n307_), .C2(new_n281_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n240_), .B2(new_n303_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT19), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n221_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n213_), .A2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n220_), .B2(new_n228_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n239_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n332_), .B(new_n335_), .C1(new_n303_), .C2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT89), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT90), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n331_), .B1(new_n303_), .B2(new_n343_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n293_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n290_), .B1(new_n355_), .B2(new_n282_), .ZN(new_n356_));
  INV_X1    g155(.A(G218gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G211gat), .ZN(new_n358_));
  INV_X1    g157(.A(G211gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G218gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n356_), .A2(new_n362_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n234_), .A2(new_n363_), .A3(new_n239_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n354_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n353_), .B1(new_n365_), .B2(new_n334_), .ZN(new_n366_));
  AOI211_X1 g165(.A(KEYINPUT87), .B(new_n335_), .C1(new_n354_), .C2(new_n364_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n344_), .B(new_n352_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT91), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n234_), .A2(new_n363_), .A3(new_n239_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n237_), .A2(new_n235_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n238_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n341_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n231_), .A2(new_n232_), .B1(new_n221_), .B2(new_n336_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n230_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n376_), .B2(new_n363_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n334_), .B1(new_n371_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT87), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n353_), .A3(new_n334_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(KEYINPUT91), .A3(new_n344_), .A4(new_n352_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n344_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n352_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n370_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n370_), .A2(new_n382_), .A3(new_n385_), .A4(KEYINPUT92), .ZN(new_n389_));
  XOR2_X1   g188(.A(G127gat), .B(G134gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(new_n247_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n278_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n263_), .A2(new_n264_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n248_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT94), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n392_), .A2(new_n395_), .A3(new_n398_), .A4(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT93), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(KEYINPUT4), .A3(new_n395_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n393_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n394_), .A2(new_n248_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n400_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT33), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n400_), .A2(new_n414_), .A3(new_n405_), .A4(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n278_), .A2(new_n391_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n408_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n392_), .A2(KEYINPUT95), .A3(new_n395_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n407_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n405_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT96), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n406_), .A2(new_n410_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n393_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n388_), .A2(new_n389_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n400_), .A2(new_n411_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n422_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n412_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n365_), .A2(new_n334_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n305_), .A2(new_n376_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n332_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n334_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n435_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n381_), .A2(new_n344_), .A3(new_n436_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n330_), .B1(new_n432_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT27), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n386_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n435_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT27), .B(new_n368_), .C1(new_n440_), .C2(new_n352_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(new_n330_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n255_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT97), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n450_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(new_n330_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n255_), .A2(new_n435_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT97), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n459_), .B(new_n255_), .C1(new_n446_), .C2(new_n452_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n454_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G29gat), .B(G36gat), .Z(new_n462_));
  XOR2_X1   g261(.A(G43gat), .B(G50gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G1gat), .A2(G8gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT14), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n464_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G113gat), .B(G141gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n482_), .B(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n461_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  INV_X1    g287(.A(G85gat), .ZN(new_n489_));
  INV_X1    g288(.A(G92gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n488_), .B(new_n491_), .C1(new_n494_), .C2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  AOI21_X1  g301(.A(new_n497_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n488_), .B1(new_n491_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n498_), .A2(new_n499_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n514_));
  XOR2_X1   g313(.A(G71gat), .B(G78gat), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n511_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n511_), .A2(new_n519_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT64), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n511_), .A2(KEYINPUT67), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n510_), .A2(new_n509_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n500_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n527_), .A2(new_n530_), .A3(KEYINPUT12), .A4(new_n519_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT68), .ZN(new_n533_));
  INV_X1    g332(.A(new_n522_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n525_), .B1(new_n534_), .B2(new_n520_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n523_), .A2(new_n536_), .A3(new_n526_), .A4(new_n531_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT13), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n528_), .A2(new_n464_), .A3(new_n500_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n527_), .A2(new_n530_), .A3(new_n465_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n550_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n550_), .A2(new_n560_), .A3(new_n551_), .A4(new_n556_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(KEYINPUT71), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n563_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT37), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n570_), .A2(new_n572_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n471_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n519_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n580_), .B(new_n585_), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n579_), .A2(KEYINPUT17), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT74), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n568_), .A2(new_n569_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n573_), .B(KEYINPUT37), .C1(new_n590_), .C2(new_n571_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n576_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n487_), .A2(new_n547_), .A3(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n593_), .A2(G1gat), .A3(new_n449_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT38), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT38), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n590_), .A2(new_n571_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n461_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n546_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n486_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT98), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n547_), .A2(new_n603_), .A3(new_n486_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n602_), .A2(new_n588_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n449_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n595_), .A2(new_n596_), .A3(new_n607_), .ZN(G1324gat));
  INV_X1    g407(.A(new_n455_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n593_), .A2(G8gat), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n611_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n598_), .A2(new_n455_), .A3(new_n605_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(G8gat), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n612_), .A2(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n615_), .A2(new_n614_), .A3(G8gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n606_), .B2(new_n255_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n593_), .A2(G15gat), .A3(new_n255_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT102), .ZN(G1326gat));
  INV_X1    g429(.A(new_n330_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G22gat), .B1(new_n606_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n631_), .A2(G22gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n593_), .B2(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(new_n597_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n589_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n600_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n487_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n435_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n576_), .A2(new_n591_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n460_), .A2(new_n458_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n430_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n444_), .B1(new_n646_), .B2(new_n389_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n451_), .B1(new_n647_), .B2(new_n330_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n459_), .B1(new_n648_), .B2(new_n255_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n643_), .B(new_n644_), .C1(new_n645_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n461_), .A2(new_n652_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n644_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n602_), .A2(new_n637_), .A3(new_n604_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n602_), .A2(new_n604_), .A3(KEYINPUT103), .A4(new_n637_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n656_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n435_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n642_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n455_), .A3(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n609_), .A2(G36gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n487_), .A2(new_n639_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n669_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n675_), .B1(new_n670_), .B2(G36gat), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  AND4_X1   g481(.A1(new_n682_), .A2(new_n671_), .A3(KEYINPUT46), .A4(new_n676_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n680_), .B2(KEYINPUT46), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n679_), .A2(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1329gat));
  INV_X1    g484(.A(new_n255_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G43gat), .B1(new_n641_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT107), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n666_), .A2(G43gat), .A3(new_n686_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n641_), .B2(new_n330_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n330_), .A2(G50gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n666_), .B2(new_n695_), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n547_), .A2(new_n486_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n589_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n598_), .A2(G57gat), .A3(new_n435_), .A4(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT110), .Z(new_n701_));
  AND2_X1   g500(.A1(new_n461_), .A2(new_n601_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n644_), .A2(new_n547_), .A3(new_n637_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n449_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n701_), .A2(new_n709_), .ZN(G1332gat));
  NAND2_X1  g509(.A1(new_n598_), .A2(new_n699_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G64gat), .B1(new_n711_), .B2(new_n609_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n609_), .A2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n704_), .B2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n711_), .B2(new_n255_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n705_), .A2(new_n243_), .A3(new_n686_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n711_), .B2(new_n631_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n631_), .A2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n704_), .B2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n697_), .A2(new_n637_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n656_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n449_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n638_), .A2(new_n547_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n702_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n489_), .A3(new_n435_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1336gat));
  OAI21_X1  g531(.A(G92gat), .B1(new_n726_), .B2(new_n609_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n490_), .A3(new_n455_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n726_), .B2(new_n255_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n737_));
  INV_X1    g536(.A(new_n502_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n729_), .A2(new_n255_), .A3(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT111), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT111), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n736_), .B(new_n737_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n742_), .B(new_n743_), .Z(G1338gat));
  NAND3_X1  g543(.A1(new_n730_), .A2(new_n501_), .A3(new_n330_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G106gat), .B1(new_n726_), .B2(new_n631_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT52), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT52), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n592_), .A2(new_n751_), .A3(new_n601_), .A4(new_n547_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n576_), .A2(new_n547_), .A3(new_n591_), .A4(new_n589_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT54), .B1(new_n753_), .B2(new_n486_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n477_), .A2(new_n475_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n485_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n546_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n545_), .A2(new_n486_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n545_), .B2(new_n486_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n533_), .A2(new_n770_), .A3(new_n537_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n533_), .A2(KEYINPUT114), .A3(new_n770_), .A4(new_n537_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n523_), .A2(new_n531_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n525_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n770_), .B2(new_n532_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n542_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n769_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n542_), .A3(new_n782_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n764_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT118), .B(new_n757_), .C1(new_n786_), .C2(new_n636_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n765_), .B(new_n766_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n778_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n783_), .B1(new_n790_), .B2(new_n544_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n636_), .B1(new_n792_), .B2(new_n763_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n793_), .B2(new_n756_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT57), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n544_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n544_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n762_), .A2(new_n545_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n796_), .A2(KEYINPUT58), .A3(new_n797_), .A4(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n644_), .A3(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n787_), .A2(new_n794_), .A3(new_n795_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n588_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n755_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n456_), .A2(new_n686_), .A3(new_n435_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n486_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT59), .B1(new_n806_), .B2(new_n807_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n806_), .C2(new_n807_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n757_), .B1(new_n786_), .B2(new_n636_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n795_), .A3(new_n803_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n755_), .B1(new_n815_), .B2(new_n637_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT120), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n815_), .A2(new_n637_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n820_), .B(new_n817_), .C1(new_n821_), .C2(new_n755_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n812_), .A2(new_n813_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n486_), .A2(G113gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT121), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n809_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n547_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n808_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n827_), .ZN(new_n829_));
  AOI221_X4 g628(.A(new_n547_), .B1(new_n819_), .B2(new_n822_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n808_), .A2(new_n832_), .A3(new_n589_), .ZN(new_n833_));
  AOI221_X4 g632(.A(new_n805_), .B1(new_n819_), .B2(new_n822_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n808_), .A2(new_n836_), .A3(new_n636_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n644_), .ZN(new_n838_));
  AOI221_X4 g637(.A(new_n838_), .B1(new_n819_), .B2(new_n822_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n839_), .B2(new_n836_), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n804_), .A2(new_n805_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n755_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n686_), .A2(new_n455_), .A3(new_n631_), .A4(new_n449_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT122), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n486_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G141gat), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n267_), .B(new_n486_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1344gat));
  OAI21_X1  g651(.A(new_n600_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G148gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n268_), .B(new_n600_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1345gat));
  OAI21_X1  g655(.A(new_n589_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n858_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n589_), .B(new_n860_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1346gat));
  OR2_X1    g661(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n838_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G162gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n847_), .A2(new_n848_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n636_), .A2(new_n866_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n865_), .A2(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n457_), .A2(new_n455_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n330_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n486_), .B(new_n871_), .C1(new_n821_), .C2(new_n755_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT62), .B(new_n215_), .C1(new_n872_), .C2(KEYINPUT22), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n872_), .B2(KEYINPUT62), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  INV_X1    g674(.A(new_n871_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n816_), .A2(new_n601_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n236_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n874_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT124), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n873_), .C1(new_n874_), .C2(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n816_), .A2(new_n876_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G176gat), .B1(new_n884_), .B2(new_n600_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n806_), .A2(new_n330_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n547_), .A2(new_n216_), .A3(new_n870_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n637_), .A2(new_n870_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n805_), .A2(new_n231_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n890_), .A2(new_n205_), .B1(new_n884_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n232_), .A3(new_n636_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n816_), .A2(new_n838_), .A3(new_n876_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n209_), .B2(new_n896_), .ZN(G1351gat));
  NOR4_X1   g696(.A1(new_n609_), .A2(new_n686_), .A3(new_n631_), .A4(new_n435_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n843_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n601_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n284_), .ZN(G1352gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n547_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n293_), .ZN(G1353gat));
  INV_X1    g702(.A(new_n899_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n588_), .B1(new_n905_), .B2(new_n359_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT126), .Z(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n359_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1354gat));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n899_), .A2(new_n838_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n357_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n899_), .A2(G218gat), .A3(new_n597_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n911_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n904_), .A2(new_n357_), .A3(new_n636_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n916_), .B(KEYINPUT127), .C1(new_n357_), .C2(new_n912_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1355gat));
endmodule


