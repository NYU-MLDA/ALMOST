//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(KEYINPUT106), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT84), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n209_), .B1(new_n212_), .B2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n210_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n207_), .B(KEYINPUT85), .C1(new_n210_), .C2(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n217_), .A2(new_n218_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n219_), .B2(KEYINPUT23), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT87), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(new_n204_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n231_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n227_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G197gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT90), .B1(new_n241_), .B2(G204gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243_));
  INV_X1    g042(.A(G204gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(G204gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT21), .ZN(new_n248_));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(G197gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n246_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(KEYINPUT21), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n247_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n240_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT95), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n208_), .A2(new_n211_), .B1(new_n206_), .B2(new_n203_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT94), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n230_), .A2(new_n225_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n237_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n256_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n260_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT19), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n240_), .A2(KEYINPUT95), .A3(new_n256_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n259_), .A2(new_n268_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n264_), .A2(new_n265_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n256_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n227_), .A2(new_n239_), .A3(new_n267_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT20), .A3(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n270_), .B(KEYINPUT93), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G8gat), .B(G36gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n273_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT97), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT97), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n273_), .A2(new_n279_), .A3(new_n288_), .A4(new_n285_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n285_), .B1(new_n273_), .B2(new_n279_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI211_X1 g091(.A(KEYINPUT98), .B(new_n285_), .C1(new_n273_), .C2(new_n279_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n287_), .B(new_n289_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI22_X1  g102(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n298_), .A2(new_n299_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(KEYINPUT1), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n307_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n308_), .A2(KEYINPUT1), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n310_), .B(new_n301_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n256_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G228gat), .A3(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n256_), .B(new_n319_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(new_n314_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n326_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n326_), .B2(KEYINPUT29), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n331_));
  OAI22_X1  g130(.A1(new_n324_), .A2(new_n325_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(KEYINPUT92), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n330_), .A2(new_n331_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n323_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n318_), .A2(new_n338_), .A3(new_n320_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n322_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n332_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n278_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT20), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT104), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n259_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n270_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n285_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n286_), .A2(KEYINPUT27), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n296_), .A2(new_n343_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT105), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT99), .ZN(new_n356_));
  XOR2_X1   g155(.A(G127gat), .B(G134gat), .Z(new_n357_));
  XOR2_X1   g156(.A(G113gat), .B(G120gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n315_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n326_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n362_), .A3(KEYINPUT4), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n362_), .B2(KEYINPUT4), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n356_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT99), .A3(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n368_), .A2(new_n370_), .A3(new_n378_), .A4(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n240_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G15gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n361_), .B(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n386_), .A2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n352_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT105), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n343_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n355_), .A2(new_n381_), .A3(new_n394_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n394_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n315_), .A2(new_n359_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n366_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT102), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n363_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n402_), .B2(new_n363_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n360_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n406_), .A2(KEYINPUT101), .A3(new_n376_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT101), .B1(new_n406_), .B2(new_n376_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n404_), .A2(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT103), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT103), .ZN(new_n411_));
  OAI221_X1 g210(.A(new_n411_), .B1(new_n407_), .B2(new_n408_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n379_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n379_), .A2(new_n414_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n290_), .B(new_n291_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n287_), .A2(new_n289_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n273_), .A2(new_n423_), .A3(new_n279_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n347_), .A2(new_n349_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n380_), .B(new_n424_), .C1(new_n425_), .C2(new_n423_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n342_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n342_), .A2(new_n381_), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n428_), .B(new_n352_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n399_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n398_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G29gat), .B(G36gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n432_), .A2(KEYINPUT76), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(KEYINPUT76), .ZN(new_n434_));
  XOR2_X1   g233(.A(G43gat), .B(G50gat), .Z(new_n435_));
  OR3_X1    g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT15), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G22gat), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  INV_X1    g240(.A(G8gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT14), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G8gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n436_), .A2(new_n437_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT15), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT81), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n438_), .A2(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G229gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n447_), .B(new_n446_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n451_), .A2(new_n455_), .B1(new_n457_), .B2(new_n454_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  OR2_X1    g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n451_), .A2(new_n455_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n454_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n461_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(KEYINPUT82), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n462_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n202_), .B1(new_n431_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  AOI211_X1 g270(.A(KEYINPUT106), .B(new_n471_), .C1(new_n398_), .C2(new_n430_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  OR3_X1    g273(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n475_), .B(new_n476_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n474_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n474_), .A3(new_n485_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n481_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n479_), .B(KEYINPUT6), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(KEYINPUT65), .A3(new_n476_), .A4(new_n475_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n492_), .A2(KEYINPUT66), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT66), .B1(new_n492_), .B2(new_n494_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT9), .B1(new_n482_), .B2(new_n483_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n486_), .B2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n498_), .A2(new_n493_), .A3(new_n501_), .A4(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT70), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n497_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n439_), .A3(new_n449_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n481_), .A2(new_n491_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n490_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n494_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n492_), .A2(KEYINPUT66), .A3(new_n494_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n488_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n505_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n447_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n508_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT77), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n518_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n508_), .A2(new_n518_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT77), .B1(new_n517_), .B2(new_n447_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(new_n529_), .B2(new_n523_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n531_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n531_), .A2(KEYINPUT78), .A3(new_n535_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT78), .B1(new_n531_), .B2(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n537_), .B(new_n541_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G57gat), .ZN(new_n547_));
  INV_X1    g346(.A(G57gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G64gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n549_), .A3(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT68), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT11), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT11), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n548_), .A2(G64gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n546_), .A2(G57gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G71gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(G78gat), .ZN(new_n562_));
  INV_X1    g361(.A(G78gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G71gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n556_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT11), .B1(new_n547_), .B2(new_n549_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n567_), .A2(KEYINPUT67), .A3(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n555_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT67), .B1(new_n567_), .B2(new_n568_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n565_), .B(new_n556_), .C1(new_n552_), .C2(KEYINPUT11), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(new_n551_), .A3(new_n554_), .A4(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(KEYINPUT69), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT69), .B1(new_n570_), .B2(new_n573_), .ZN(new_n576_));
  NOR4_X1   g375(.A1(new_n515_), .A2(new_n575_), .A3(new_n576_), .A4(new_n516_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n505_), .B(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n515_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n582_));
  INV_X1    g381(.A(new_n573_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n571_), .A2(new_n572_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n570_), .A2(KEYINPUT71), .A3(new_n573_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT12), .A3(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n578_), .B1(new_n581_), .B2(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n570_), .A2(KEYINPUT71), .A3(new_n573_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT71), .B1(new_n570_), .B2(new_n573_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n507_), .A3(KEYINPUT72), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n577_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT69), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n497_), .A2(new_n505_), .B1(new_n596_), .B2(new_n574_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT73), .B1(new_n597_), .B2(KEYINPUT12), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n515_), .A2(new_n516_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n591_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n577_), .B2(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G120gat), .B(G148gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(new_n606_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(KEYINPUT13), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n589_), .A2(new_n590_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n446_), .B(new_n628_), .Z(new_n629_));
  AOI211_X1 g428(.A(new_n621_), .B(new_n626_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n575_), .A2(new_n576_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n629_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n545_), .A2(new_n620_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n473_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n441_), .A3(new_n380_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n540_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n398_), .B2(new_n430_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT107), .B1(new_n620_), .B2(new_n471_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n637_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n618_), .A2(new_n648_), .A3(new_n469_), .A4(new_n619_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n645_), .A2(KEYINPUT108), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT108), .B1(new_n645_), .B2(new_n650_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n380_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G1gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n641_), .A2(new_n642_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n643_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(new_n395_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n442_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n645_), .A2(new_n657_), .A3(new_n650_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G8gat), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n659_), .A3(G8gat), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n639_), .A2(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g463(.A1(new_n640_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n394_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(G15gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT41), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT41), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(new_n342_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G22gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G22gat), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n343_), .A2(G22gat), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n673_), .A2(new_n674_), .B1(new_n639_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI221_X1 g477(.A(KEYINPUT109), .B1(new_n639_), .B2(new_n675_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n646_), .A2(new_n637_), .A3(new_n649_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n431_), .B2(new_n545_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n543_), .A2(new_n544_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT43), .B(new_n685_), .C1(new_n398_), .C2(new_n430_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n682_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n380_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n644_), .A2(new_n637_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n620_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n381_), .A2(G29gat), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n694_), .B(new_n695_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n681_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n696_), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT110), .B(new_n698_), .C1(new_n691_), .C2(G29gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n657_), .A3(new_n690_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n395_), .A2(G36gat), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n694_), .B(new_n703_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n473_), .A2(new_n694_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n399_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n689_), .A2(G43gat), .A3(new_n394_), .A4(new_n690_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n712_), .B2(new_n343_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n689_), .A2(G50gat), .A3(new_n342_), .A4(new_n690_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  INV_X1    g520(.A(new_n620_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n469_), .A3(new_n637_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n645_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT112), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n645_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n380_), .A2(G57gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n721_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n545_), .A2(new_n637_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n620_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n469_), .B1(new_n398_), .B2(new_n430_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n548_), .B1(new_n736_), .B2(new_n381_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n728_), .A2(new_n721_), .A3(new_n729_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(new_n736_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n546_), .A3(new_n657_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n657_), .A3(new_n727_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G64gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n561_), .A3(new_n394_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n725_), .A2(new_n394_), .A3(new_n727_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G71gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n741_), .A2(new_n563_), .A3(new_n342_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n725_), .A2(new_n342_), .A3(new_n727_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G78gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT114), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n693_), .A2(new_n722_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n734_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n482_), .A3(new_n380_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n684_), .A2(new_n686_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n722_), .A2(new_n469_), .A3(new_n647_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n380_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n766_), .B1(new_n772_), .B2(new_n482_), .ZN(G1336gat));
  AOI21_X1  g572(.A(G92gat), .B1(new_n765_), .B2(new_n657_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n657_), .A2(G92gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT116), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n775_), .A2(new_n776_), .B1(new_n770_), .B2(new_n778_), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n769_), .B2(new_n399_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n765_), .A2(new_n394_), .A3(new_n502_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(G1338gat));
  OAI211_X1 g583(.A(new_n342_), .B(new_n768_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G106gat), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n734_), .A2(new_n503_), .A3(new_n342_), .A4(new_n764_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT118), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g592(.A1(new_n685_), .A2(new_n471_), .A3(new_n722_), .A4(new_n647_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n638_), .A2(new_n471_), .A3(new_n795_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n461_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n456_), .B2(new_n454_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT122), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n452_), .A2(new_n453_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n451_), .A2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n465_), .A2(KEYINPUT82), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n458_), .A2(new_n467_), .A3(new_n461_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n616_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n597_), .A2(KEYINPUT73), .A3(KEYINPUT12), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n600_), .B1(new_n599_), .B2(new_n591_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n517_), .A2(new_n632_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n581_), .A2(new_n587_), .A3(new_n578_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT72), .B1(new_n592_), .B2(new_n507_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n605_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n604_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n594_), .A2(new_n602_), .A3(KEYINPUT55), .A4(new_n603_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n594_), .A2(new_n602_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT120), .A3(new_n605_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n612_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n469_), .A2(new_n615_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n825_), .B2(new_n612_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT56), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n809_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n540_), .B1(KEYINPUT124), .B2(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n809_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n828_), .B1(new_n832_), .B2(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT120), .B1(new_n823_), .B2(new_n605_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n818_), .B(new_n603_), .C1(new_n594_), .C2(new_n602_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n821_), .A2(new_n822_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n614_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n849_), .B2(new_n831_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n842_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n841_), .B1(new_n851_), .B2(new_n835_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n825_), .A2(new_n844_), .A3(new_n612_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n808_), .A2(new_n615_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n853_), .A2(KEYINPUT58), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n808_), .A2(new_n615_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n849_), .B2(new_n844_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(KEYINPUT58), .A4(new_n853_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n854_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n849_), .A2(new_n844_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n857_), .A2(new_n545_), .A3(new_n861_), .A4(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n840_), .A2(new_n852_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n799_), .B1(new_n867_), .B2(new_n637_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n381_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n355_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .A4(new_n469_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n637_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n799_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n380_), .A3(new_n871_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n869_), .A2(KEYINPUT59), .A3(new_n871_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n471_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n872_), .B1(new_n880_), .B2(new_n870_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n882_), .A2(KEYINPUT60), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n722_), .B2(KEYINPUT60), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n869_), .A2(new_n871_), .A3(new_n883_), .A4(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n722_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n869_), .A2(new_n888_), .A3(new_n871_), .A4(new_n647_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n637_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n888_), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n869_), .A2(new_n892_), .A3(new_n871_), .A4(new_n644_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n685_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n892_), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n657_), .A2(new_n343_), .A3(new_n394_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n869_), .A2(new_n469_), .A3(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n869_), .A2(new_n620_), .A3(new_n896_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n869_), .A2(new_n647_), .A3(new_n896_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  NAND2_X1  g702(.A1(new_n869_), .A2(new_n896_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G162gat), .B1(new_n904_), .B2(new_n685_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n540_), .A2(G162gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(new_n906_), .ZN(G1347gat));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n395_), .A2(new_n399_), .A3(new_n342_), .A4(new_n380_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n875_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n471_), .ZN(new_n911_));
  INV_X1    g710(.A(G169gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n908_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n234_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(G169gat), .C1(new_n910_), .C2(new_n471_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  NOR2_X1   g715(.A1(new_n910_), .A2(new_n722_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n918_));
  OR2_X1    g717(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  INV_X1    g720(.A(new_n909_), .ZN(new_n922_));
  NOR4_X1   g721(.A1(new_n868_), .A2(new_n211_), .A3(new_n637_), .A4(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n910_), .A2(new_n637_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n924_), .B(new_n925_), .C1(new_n926_), .C2(G183gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n868_), .A2(new_n922_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G183gat), .B1(new_n928_), .B2(new_n647_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT126), .B1(new_n929_), .B2(new_n923_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n910_), .B2(new_n685_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n208_), .A3(new_n644_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1351gat));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n395_), .A2(new_n428_), .A3(new_n394_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n875_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n868_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940_), .B2(new_n469_), .ZN(new_n941_));
  AOI211_X1 g740(.A(new_n241_), .B(new_n471_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1352gat));
  AOI21_X1  g742(.A(new_n935_), .B1(new_n875_), .B2(new_n936_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n868_), .A2(KEYINPUT127), .A3(new_n938_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G204gat), .B1(new_n946_), .B2(new_n722_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n940_), .A2(new_n244_), .A3(new_n620_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1353gat));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n637_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n940_), .B2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n952_), .ZN(new_n954_));
  AOI211_X1 g753(.A(new_n950_), .B(new_n954_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n946_), .B2(new_n685_), .ZN(new_n957_));
  INV_X1    g756(.A(G218gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n940_), .A2(new_n958_), .A3(new_n644_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n959_), .ZN(G1355gat));
endmodule


