//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT35), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  INV_X1    g008(.A(G43gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G50gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n209_), .B(G43gat), .ZN(new_n213_));
  INV_X1    g012(.A(G50gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n215_), .A3(KEYINPUT15), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G85gat), .B(G92gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n231_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(new_n232_), .C2(KEYINPUT9), .ZN(new_n238_));
  AND3_X1   g037(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT10), .B(G99gat), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n241_), .B(new_n242_), .C1(G106gat), .C2(new_n243_), .ZN(new_n244_));
  OAI22_X1  g043(.A1(new_n234_), .A2(new_n235_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n208_), .B1(new_n220_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n216_), .A2(new_n245_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n230_), .A2(new_n233_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n237_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT9), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT64), .B(new_n252_), .C1(new_n233_), .C2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n222_), .A2(KEYINPUT10), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT10), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G99gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(G106gat), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n227_), .A2(new_n228_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n242_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n250_), .A2(new_n251_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  AOI211_X1 g061(.A(KEYINPUT70), .B(new_n262_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n202_), .B(new_n207_), .C1(new_n248_), .C2(new_n263_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n246_), .A2(new_n263_), .A3(new_n247_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n207_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n220_), .A2(new_n245_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n247_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n205_), .A2(new_n206_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n207_), .B(KEYINPUT72), .Z(new_n271_));
  NAND4_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G190gat), .B(G218gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G134gat), .ZN(new_n275_));
  INV_X1    g074(.A(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT74), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n264_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n277_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT36), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n280_), .A2(KEYINPUT75), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n273_), .A2(new_n285_), .A3(new_n279_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT37), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n264_), .A2(new_n267_), .A3(new_n272_), .A4(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n280_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n281_), .A2(KEYINPUT73), .A3(new_n283_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G15gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT77), .B(G1gat), .Z(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(G57gat), .ZN(new_n305_));
  INV_X1    g104(.A(G64gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G57gat), .A2(G64gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n311_));
  INV_X1    g110(.A(G71gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G78gat), .ZN(new_n313_));
  INV_X1    g112(.A(G78gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G71gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n310_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n310_), .B2(new_n316_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n309_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G57gat), .A2(G64gat), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT11), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G71gat), .B(G78gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT65), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n310_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n319_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n304_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT16), .B(G183gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G211gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(G127gat), .B(G155gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n332_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n332_), .A2(new_n338_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT78), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n294_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT79), .ZN(new_n345_));
  XOR2_X1   g144(.A(G15gat), .B(G43gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT23), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(KEYINPUT23), .ZN(new_n353_));
  MUX2_X1   g152(.A(new_n352_), .B(new_n353_), .S(KEYINPUT82), .Z(new_n354_));
  INV_X1    g153(.A(G169gat), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT24), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT81), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(G190gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT25), .B(G183gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G190gat), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n365_), .B(new_n366_), .C1(new_n367_), .C2(new_n363_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n360_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n354_), .A2(new_n362_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n353_), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n359_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G169gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n356_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT83), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n378_), .A2(new_n380_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n387_), .B2(new_n386_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT31), .Z(new_n391_));
  NOR3_X1   g190(.A1(new_n382_), .A2(new_n383_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n377_), .B(KEYINPUT83), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n379_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n395_), .B2(new_n381_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n350_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n391_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n381_), .A3(new_n393_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n349_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G141gat), .ZN(new_n403_));
  INV_X1    g202(.A(G148gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT86), .B1(new_n405_), .B2(KEYINPUT85), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n405_), .B2(KEYINPUT86), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(KEYINPUT2), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(KEYINPUT2), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n410_), .A2(new_n411_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n412_));
  OAI211_X1 g211(.A(G141gat), .B(G148gat), .C1(new_n409_), .C2(KEYINPUT2), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT86), .B(KEYINPUT3), .C1(new_n405_), .C2(KEYINPUT85), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n408_), .A2(new_n412_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT1), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n416_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n405_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT29), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G22gat), .B(G50gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n426_), .B(KEYINPUT28), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n425_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT21), .ZN(new_n431_));
  XOR2_X1   g230(.A(G197gat), .B(G204gat), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n431_), .A2(new_n432_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n424_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G228gat), .A3(G233gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G228gat), .A2(G233gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n440_), .B(new_n435_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G78gat), .B(G106gat), .Z(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(KEYINPUT89), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n428_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n443_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT88), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n428_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n439_), .A2(new_n441_), .A3(new_n451_), .A4(new_n443_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n366_), .A2(new_n367_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n456_), .A2(new_n353_), .A3(new_n358_), .A4(new_n360_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT90), .Z(new_n458_));
  OAI21_X1  g257(.A(new_n354_), .B1(G183gat), .B2(G190gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n375_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n435_), .ZN(new_n462_));
  OAI211_X1 g261(.A(KEYINPUT20), .B(new_n462_), .C1(new_n378_), .C2(new_n435_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT20), .B1(new_n461_), .B2(new_n435_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n378_), .A2(new_n435_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT18), .B(G64gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G92gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G8gat), .B(G36gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT0), .B(G57gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G85gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G29gat), .Z(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n424_), .A2(new_n484_), .A3(new_n390_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n424_), .A2(new_n390_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT91), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n386_), .A2(new_n388_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n436_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n424_), .A2(new_n494_), .A3(new_n390_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT4), .A4(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n483_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n495_), .A3(new_n493_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(new_n483_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT33), .B(new_n482_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n466_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n477_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n496_), .A2(new_n488_), .A3(new_n487_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n483_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n504_), .B1(new_n507_), .B2(new_n481_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n498_), .A2(new_n483_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(new_n481_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n512_));
  OAI211_X1 g311(.A(KEYINPUT94), .B(new_n504_), .C1(new_n507_), .C2(new_n481_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n502_), .A2(new_n510_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n507_), .B(new_n481_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n475_), .A2(KEYINPUT32), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n460_), .A2(new_n457_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n469_), .B(KEYINPUT20), .C1(new_n435_), .C2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n519_), .A2(new_n465_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n463_), .A2(new_n465_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n515_), .B(new_n522_), .C1(new_n471_), .C2(new_n517_), .ZN(new_n523_));
  AOI211_X1 g322(.A(new_n402_), .B(new_n455_), .C1(new_n514_), .C2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n401_), .B(new_n454_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n476_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(KEYINPUT27), .A3(new_n501_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n477_), .A2(new_n501_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT27), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n525_), .A2(new_n531_), .A3(new_n515_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n304_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n303_), .B(new_n299_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n220_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n216_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n355_), .ZN(new_n544_));
  INV_X1    g343(.A(G197gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n542_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n250_), .A2(new_n251_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n254_), .A2(new_n261_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n320_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n326_), .A2(new_n327_), .A3(new_n319_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT66), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n329_), .A2(new_n555_), .A3(new_n262_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n245_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT67), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT12), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n245_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n561_), .C1(new_n558_), .C2(new_n245_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n560_), .A2(new_n561_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n356_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n548_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n533_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n345_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n515_), .A3(new_n298_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n284_), .A2(new_n286_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n284_), .A2(KEYINPUT96), .A3(new_n286_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n342_), .ZN(new_n598_));
  NOR4_X1   g397(.A1(new_n533_), .A2(new_n597_), .A3(new_n587_), .A4(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n302_), .B1(new_n599_), .B2(new_n515_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n592_), .A2(new_n600_), .ZN(G1324gat));
  NAND3_X1  g400(.A1(new_n589_), .A2(new_n299_), .A3(new_n531_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT97), .Z(new_n603_));
  AOI21_X1  g402(.A(new_n299_), .B1(new_n599_), .B2(new_n531_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT39), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(G1325gat));
  AOI21_X1  g407(.A(new_n296_), .B1(new_n599_), .B2(new_n402_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT98), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT41), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n589_), .A2(new_n296_), .A3(new_n402_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n454_), .B(KEYINPUT99), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n599_), .B2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT42), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n589_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1327gat));
  AOI21_X1  g418(.A(new_n343_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n588_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G29gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n515_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n287_), .A2(new_n293_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n624_), .B(new_n625_), .C1(new_n524_), .C2(new_n532_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT100), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT43), .B1(new_n533_), .B2(new_n294_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n531_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n515_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n402_), .A2(new_n454_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n455_), .A2(new_n401_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n629_), .B(new_n630_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n514_), .A2(new_n523_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n401_), .A3(new_n454_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n625_), .A4(new_n624_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n627_), .A2(new_n628_), .A3(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n587_), .A2(new_n343_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n640_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n515_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n645_), .B2(G29gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n623_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n531_), .B(KEYINPUT103), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n621_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT45), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n531_), .A3(new_n644_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(G36gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n654_), .B2(G36gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT46), .B(new_n653_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1329gat));
  NAND4_X1  g461(.A1(new_n643_), .A2(G43gat), .A3(new_n402_), .A4(new_n644_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n621_), .A2(new_n402_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n210_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT104), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n668_), .A3(new_n665_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(KEYINPUT47), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT47), .B1(new_n667_), .B2(new_n669_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1330gat));
  AOI21_X1  g471(.A(G50gat), .B1(new_n621_), .B2(new_n615_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n643_), .A2(G50gat), .A3(new_n644_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n455_), .ZN(G1331gat));
  NOR2_X1   g474(.A1(new_n533_), .A2(new_n597_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n586_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n547_), .A3(new_n677_), .A4(new_n343_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(new_n305_), .A3(new_n630_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n636_), .A2(new_n547_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT105), .Z(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n586_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n345_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(KEYINPUT106), .A3(new_n345_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n515_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n687_), .B2(new_n305_), .ZN(G1332gat));
  INV_X1    g487(.A(new_n651_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G64gat), .B1(new_n678_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n686_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n651_), .A2(new_n306_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(G1333gat));
  OAI21_X1  g493(.A(G71gat), .B1(new_n678_), .B2(new_n401_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT49), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n402_), .A2(new_n312_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n692_), .B2(new_n697_), .ZN(G1334gat));
  INV_X1    g497(.A(new_n615_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G78gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n685_), .A2(new_n686_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G78gat), .B1(new_n678_), .B2(new_n699_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(KEYINPUT107), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1335gat));
  NAND2_X1  g507(.A1(new_n682_), .A2(new_n620_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n709_), .A2(G85gat), .A3(new_n630_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  INV_X1    g510(.A(new_n343_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n548_), .A2(new_n586_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n639_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n515_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G85gat), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n710_), .A2(new_n711_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n711_), .B1(new_n710_), .B2(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1336gat));
  INV_X1    g518(.A(new_n709_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G92gat), .B1(new_n720_), .B2(new_n531_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n714_), .A2(G92gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n651_), .B2(new_n722_), .ZN(G1337gat));
  NOR2_X1   g522(.A1(new_n401_), .A2(new_n243_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n714_), .A2(new_n402_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G99gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT109), .B(new_n222_), .C1(new_n714_), .C2(new_n402_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n725_), .B(new_n732_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n720_), .A2(new_n223_), .A3(new_n455_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n639_), .A2(new_n455_), .A3(new_n712_), .A4(new_n713_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n736_), .B(G106gat), .C1(KEYINPUT110), .C2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n737_), .A2(KEYINPUT110), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n735_), .A2(new_n740_), .A3(new_n744_), .A4(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT59), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n629_), .A2(new_n515_), .A3(new_n632_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT118), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n558_), .A2(new_n245_), .A3(new_n565_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n558_), .A2(new_n245_), .B1(new_n562_), .B2(KEYINPUT12), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n752_), .B(new_n561_), .C1(new_n755_), .C2(new_n557_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n555_), .B1(new_n329_), .B2(new_n262_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n558_), .A2(new_n245_), .A3(KEYINPUT66), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n566_), .B(new_n564_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n561_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT111), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n572_), .B2(new_n567_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n561_), .B1(new_n558_), .B2(new_n245_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT68), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n569_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n755_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n751_), .B1(new_n762_), .B2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n757_), .A2(new_n758_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n760_), .B1(new_n771_), .B2(new_n567_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n752_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n759_), .A2(KEYINPUT111), .A3(new_n760_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n755_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT55), .B1(new_n767_), .B2(new_n755_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n778_), .A3(KEYINPUT112), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n578_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT113), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n770_), .A2(new_n779_), .A3(KEYINPUT56), .A4(new_n578_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n762_), .A2(new_n769_), .A3(new_n751_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT112), .B1(new_n775_), .B2(new_n778_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n578_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n780_), .A2(new_n791_), .A3(new_n781_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n783_), .A2(new_n786_), .A3(new_n790_), .A4(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n548_), .A3(new_n580_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n541_), .A2(new_n537_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n534_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n546_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n546_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n542_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n582_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n597_), .B1(new_n794_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n782_), .A2(new_n784_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n802_), .A2(KEYINPUT58), .A3(new_n580_), .A4(new_n799_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n579_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n799_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT58), .B1(new_n806_), .B2(new_n799_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n294_), .A2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(KEYINPUT57), .A2(new_n801_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n800_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n780_), .A2(new_n791_), .A3(new_n781_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n791_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n784_), .B(KEYINPUT114), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n547_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n814_), .B1(new_n819_), .B2(new_n580_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n813_), .B1(new_n820_), .B2(new_n597_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n343_), .B1(new_n811_), .B2(new_n821_), .ZN(new_n822_));
  AND4_X1   g621(.A1(new_n547_), .A2(new_n294_), .A3(new_n586_), .A4(new_n343_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT54), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n748_), .B(new_n750_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n801_), .B2(new_n812_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT116), .B(new_n813_), .C1(new_n820_), .C2(new_n597_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n811_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n598_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n824_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n749_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n548_), .B(new_n825_), .C1(new_n832_), .C2(new_n748_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G113gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n824_), .B1(new_n829_), .B2(new_n598_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n835_), .A2(G113gat), .A3(new_n547_), .A4(new_n749_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n747_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT119), .B(new_n836_), .C1(new_n833_), .C2(G113gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n832_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n835_), .B2(new_n749_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n844_), .A2(new_n677_), .A3(new_n825_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n832_), .B2(new_n343_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT120), .B(G127gat), .Z(new_n848_));
  AND3_X1   g647(.A1(new_n844_), .A2(new_n825_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n342_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n832_), .B2(new_n597_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n844_), .A2(new_n624_), .A3(new_n825_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g652(.A(new_n631_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n835_), .A2(new_n630_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n689_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n547_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT121), .B(G141gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n586_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT122), .B(G148gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n856_), .A2(new_n712_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT123), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n863_), .B(new_n865_), .ZN(G1346gat));
  NOR3_X1   g665(.A1(new_n856_), .A2(new_n276_), .A3(new_n294_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n855_), .A2(new_n597_), .A3(new_n689_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n276_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n689_), .A2(new_n515_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n402_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n699_), .B(new_n873_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n547_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n870_), .B1(new_n875_), .B2(new_n355_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n374_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT62), .B(G169gat), .C1(new_n874_), .C2(new_n547_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  INV_X1    g678(.A(new_n874_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G176gat), .B1(new_n880_), .B2(new_n677_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n835_), .A2(new_n455_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n872_), .A2(new_n356_), .A3(new_n586_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  OR3_X1    g683(.A1(new_n874_), .A2(new_n366_), .A3(new_n598_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n885_), .A2(KEYINPUT124), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(KEYINPUT124), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n872_), .A2(new_n712_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G183gat), .B1(new_n882_), .B2(new_n888_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n886_), .A2(new_n887_), .A3(new_n889_), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n874_), .B2(new_n294_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n597_), .A2(new_n367_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n874_), .B2(new_n892_), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n835_), .A2(new_n854_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n894_), .A2(new_n548_), .A3(new_n871_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(new_n545_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT125), .B(G197gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n895_), .B2(new_n898_), .ZN(G1352gat));
  AND2_X1   g698(.A1(new_n894_), .A2(new_n871_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n677_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n830_), .A2(new_n831_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n598_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n904_), .A2(new_n631_), .A3(new_n871_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT126), .ZN(new_n907_));
  INV_X1    g706(.A(G211gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n894_), .A2(new_n909_), .A3(new_n871_), .A4(new_n905_), .ZN(new_n910_));
  AND4_X1   g709(.A1(new_n903_), .A2(new_n907_), .A3(new_n908_), .A4(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n907_), .A2(new_n910_), .B1(new_n903_), .B2(new_n908_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1354gat));
  AOI21_X1  g712(.A(G218gat), .B1(new_n900_), .B2(new_n597_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n624_), .A2(G218gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT127), .Z(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n900_), .B2(new_n916_), .ZN(G1355gat));
endmodule


