//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT91), .B(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G197gat), .B2(G204gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n205_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n206_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(G204gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n211_), .B1(new_n214_), .B2(KEYINPUT21), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT82), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n224_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n230_), .B(KEYINPUT81), .ZN(new_n234_));
  INV_X1    g033(.A(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(G176gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(KEYINPUT97), .B2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(KEYINPUT97), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n233_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT26), .B(G190gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT96), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT25), .B(G183gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n221_), .A2(new_n228_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n204_), .B1(new_n219_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT101), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n217_), .B(KEYINPUT92), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT80), .B(G190gat), .Z(new_n250_));
  OAI21_X1  g049(.A(new_n229_), .B1(new_n250_), .B2(G183gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n221_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n234_), .A2(new_n231_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n227_), .B(new_n253_), .C1(new_n234_), .C2(new_n237_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n222_), .A2(KEYINPUT25), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT79), .Z(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n250_), .B2(KEYINPUT26), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n222_), .A2(KEYINPUT25), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n249_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n246_), .A2(new_n247_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n203_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n217_), .ZN(new_n266_));
  OAI221_X1 g065(.A(KEYINPUT20), .B1(new_n266_), .B2(new_n245_), .C1(new_n249_), .C2(new_n261_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(new_n203_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT18), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n204_), .B(new_n203_), .C1(new_n245_), .C2(new_n266_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n262_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT99), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT98), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n267_), .A2(new_n280_), .A3(new_n203_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n249_), .A2(new_n261_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT20), .B1(new_n245_), .B2(new_n266_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n203_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT98), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n279_), .A2(new_n273_), .A3(new_n281_), .A4(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n275_), .A2(KEYINPUT27), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n277_), .B(KEYINPUT99), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n281_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n274_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n286_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT102), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT102), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n294_), .B(KEYINPUT27), .C1(new_n290_), .C2(new_n286_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n287_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n300_), .B(new_n301_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(KEYINPUT85), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT88), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n308_), .A2(KEYINPUT86), .A3(KEYINPUT1), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT86), .B1(new_n308_), .B2(KEYINPUT1), .ZN(new_n312_));
  OAI221_X1 g111(.A(new_n309_), .B1(KEYINPUT1), .B2(new_n308_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(new_n305_), .C1(G141gat), .C2(G148gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT87), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT84), .B1(new_n317_), .B2(new_n318_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n310_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n324_), .A2(KEYINPUT4), .A3(new_n326_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT100), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n324_), .A2(KEYINPUT100), .A3(KEYINPUT4), .A4(new_n326_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n336_), .B2(new_n329_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n337_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n323_), .B(KEYINPUT31), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(KEYINPUT83), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G15gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT30), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n345_), .B(new_n349_), .Z(new_n350_));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n261_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n350_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n357_));
  INV_X1    g156(.A(new_n219_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G233gat), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(KEYINPUT90), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(KEYINPUT90), .ZN(new_n362_));
  OAI21_X1  g161(.A(G228gat), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n249_), .A2(new_n363_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n359_), .A2(new_n364_), .B1(new_n357_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n368_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(KEYINPUT94), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n316_), .B2(KEYINPUT29), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n310_), .A2(new_n315_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n376_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n374_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT94), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n366_), .A2(new_n386_), .A3(new_n368_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n366_), .A2(new_n389_), .A3(new_n368_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n389_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n370_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(new_n385_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n372_), .A2(new_n388_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n296_), .A2(new_n356_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n336_), .A2(new_n328_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n325_), .A2(new_n327_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n341_), .B1(new_n398_), .B2(new_n329_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT33), .B1(new_n337_), .B2(new_n341_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n337_), .A2(KEYINPUT33), .A3(new_n341_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n337_), .B(new_n341_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n273_), .A2(KEYINPUT32), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n288_), .A2(new_n289_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n403_), .A2(new_n404_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n395_), .A2(new_n343_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n410_), .A2(new_n395_), .B1(new_n296_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n355_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n396_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT72), .B(G15gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G22gat), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G1gat), .B(G8gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G29gat), .B(G36gat), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n425_), .A2(KEYINPUT70), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(KEYINPUT70), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G43gat), .B(G50gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n424_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n424_), .A2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n416_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n422_), .B(new_n423_), .Z(new_n437_));
  INV_X1    g236(.A(KEYINPUT15), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n425_), .B(KEYINPUT70), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(KEYINPUT15), .A3(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n415_), .A3(new_n433_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n446_), .A3(KEYINPUT78), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n445_), .A2(new_n448_), .A3(new_n433_), .A4(new_n415_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G141gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G169gat), .B(G197gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n449_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT64), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT64), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n470_));
  INV_X1    g269(.A(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G85gat), .ZN(new_n474_));
  INV_X1    g273(.A(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT9), .A3(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n459_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT64), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT64), .B1(new_n466_), .B2(new_n467_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n473_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n488_));
  INV_X1    g287(.A(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n471_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n465_), .A2(new_n492_), .A3(new_n468_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n476_), .A2(new_n477_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT8), .ZN(new_n495_));
  INV_X1    g294(.A(new_n494_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n462_), .A2(new_n464_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n491_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n493_), .A2(new_n495_), .B1(new_n499_), .B2(KEYINPUT8), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n487_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n432_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n495_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n484_), .B2(new_n492_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n490_), .B(new_n491_), .C1(new_n462_), .C2(new_n464_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n496_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n481_), .B(new_n486_), .C1(new_n504_), .C2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n430_), .A2(new_n438_), .A3(new_n431_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT15), .B1(new_n442_), .B2(new_n429_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n502_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n444_), .A2(new_n508_), .B1(new_n515_), .B2(new_n514_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n502_), .ZN(new_n521_));
  OAI22_X1  g320(.A1(new_n518_), .A2(new_n521_), .B1(new_n515_), .B2(new_n514_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(KEYINPUT69), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n519_), .A3(new_n502_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT35), .A4(new_n513_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G190gat), .B(G218gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(KEYINPUT36), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n533_), .ZN(new_n536_));
  AOI211_X1 g335(.A(KEYINPUT71), .B(new_n536_), .C1(new_n522_), .C2(new_n525_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n532_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT37), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n541_), .B1(new_n501_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(new_n548_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n550_), .B(new_n551_), .C1(new_n487_), .C2(new_n500_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n508_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n487_), .B2(new_n500_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n493_), .A2(new_n495_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n559_), .A2(new_n481_), .A3(new_n486_), .A4(new_n548_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(KEYINPUT66), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT66), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n501_), .A2(new_n562_), .A3(new_n548_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n541_), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n555_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n570_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT67), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(KEYINPUT67), .A3(new_n570_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT68), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT13), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n548_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT73), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n424_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT75), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  AND2_X1   g390(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n585_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n585_), .A2(new_n592_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT76), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(KEYINPUT76), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n594_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n532_), .B(new_n599_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n539_), .A2(new_n581_), .A3(new_n598_), .A4(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT77), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n414_), .A2(new_n458_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n419_), .A3(new_n405_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT38), .ZN(new_n605_));
  INV_X1    g404(.A(new_n581_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n458_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n538_), .B(KEYINPUT103), .Z(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n414_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n296_), .A2(new_n411_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n405_), .A2(new_n409_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n337_), .A2(new_n341_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n290_), .A2(new_n286_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n404_), .A4(new_n400_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n395_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n413_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n396_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n610_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT104), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n608_), .B1(new_n611_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n343_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n605_), .A2(new_n627_), .ZN(G1324gat));
  NAND3_X1  g427(.A1(new_n603_), .A2(new_n420_), .A3(new_n296_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n296_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(G8gat), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT39), .B(new_n420_), .C1(new_n625_), .C2(new_n296_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g434(.A1(new_n603_), .A2(new_n347_), .A3(new_n355_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G15gat), .B1(new_n626_), .B2(new_n413_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n603_), .A2(new_n642_), .A3(new_n395_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n392_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n388_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n644_), .A2(new_n393_), .B1(new_n645_), .B2(new_n371_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G22gat), .B1(new_n626_), .B2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n643_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  NAND2_X1  g449(.A1(new_n539_), .A2(new_n600_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n414_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(new_n411_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n287_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n294_), .B1(new_n617_), .B2(KEYINPUT27), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n291_), .A2(KEYINPUT102), .A3(new_n292_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n613_), .A2(new_n618_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n646_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n355_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n654_), .B(new_n651_), .C1(new_n663_), .C2(new_n396_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n653_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n598_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n607_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n670_), .B(new_n667_), .C1(new_n653_), .C2(new_n664_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n669_), .A2(new_n671_), .A3(new_n343_), .ZN(new_n672_));
  INV_X1    g471(.A(G29gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n538_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n606_), .A2(new_n674_), .A3(new_n598_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n622_), .A2(new_n457_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n405_), .A2(new_n673_), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n672_), .A2(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n676_), .A2(G36gat), .A3(new_n659_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT45), .Z(new_n680_));
  NAND2_X1  g479(.A1(new_n665_), .A2(new_n668_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n670_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n668_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n296_), .A4(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n669_), .A2(new_n671_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n687_), .B2(new_n296_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n680_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT46), .B(new_n680_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NAND3_X1  g492(.A1(new_n687_), .A2(G43gat), .A3(new_n355_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n676_), .A2(new_n413_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(G43gat), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g496(.A1(new_n676_), .A2(G50gat), .A3(new_n646_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n699_), .A3(new_n395_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n687_), .B2(new_n395_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1331gat));
  NAND2_X1  g502(.A1(new_n611_), .A2(new_n624_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n666_), .A2(new_n457_), .A3(new_n581_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n343_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n414_), .A2(new_n457_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n539_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n606_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n405_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n706_), .B2(new_n296_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n715_), .A3(new_n296_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n720_), .A3(new_n355_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G71gat), .B1(new_n707_), .B2(new_n413_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT49), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT49), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n726_), .A3(new_n395_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n706_), .A2(new_n395_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(G78gat), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT108), .B(new_n727_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n581_), .A2(new_n598_), .A3(new_n457_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n665_), .A2(new_n737_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT109), .Z(new_n739_));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n343_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n581_), .A2(new_n674_), .A3(new_n598_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n709_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n474_), .A3(new_n405_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n740_), .A2(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n739_), .B2(new_n659_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n475_), .A3(new_n296_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1337gat));
  AOI21_X1  g547(.A(new_n489_), .B1(new_n738_), .B2(new_n355_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n355_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n743_), .B2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g551(.A1(new_n665_), .A2(new_n395_), .A3(new_n737_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT110), .B1(new_n753_), .B2(G106gat), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT110), .A3(G106gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n742_), .A2(G106gat), .A3(new_n646_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n758_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n710_), .A2(new_n765_), .A3(new_n458_), .A4(new_n581_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT54), .B1(new_n601_), .B2(new_n457_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n415_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n445_), .A2(new_n416_), .A3(new_n433_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n455_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n454_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n569_), .A2(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n556_), .A2(KEYINPUT12), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n552_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n540_), .B1(new_n777_), .B2(new_n560_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n560_), .A2(new_n540_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n776_), .B2(new_n552_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(KEYINPUT55), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n555_), .A2(KEYINPUT112), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n549_), .B(KEYINPUT55), .C1(new_n553_), .C2(new_n554_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(KEYINPUT113), .A3(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n775_), .B1(new_n785_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n570_), .B1(new_n785_), .B2(new_n790_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n774_), .A2(new_n791_), .B1(new_n792_), .B2(KEYINPUT56), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n791_), .A2(new_n774_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n773_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n773_), .B(KEYINPUT58), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n651_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(new_n778_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n781_), .A2(new_n779_), .A3(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT112), .B1(new_n555_), .B2(new_n783_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n788_), .A2(new_n789_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n569_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n791_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n574_), .A2(new_n575_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n457_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n801_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n454_), .A2(new_n456_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n792_), .A2(KEYINPUT56), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n813_), .B(KEYINPUT114), .C1(new_n814_), .C2(new_n791_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n576_), .A2(new_n772_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n674_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n797_), .A2(new_n822_), .A3(new_n651_), .A4(new_n798_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n800_), .A2(new_n820_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n768_), .B1(new_n824_), .B2(new_n666_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n659_), .A2(new_n405_), .A3(new_n646_), .A4(new_n355_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n457_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT117), .Z(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n826_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n825_), .C2(new_n826_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n820_), .A2(new_n821_), .A3(new_n799_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n768_), .B1(new_n835_), .B2(new_n666_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n842_), .A3(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n457_), .A2(G113gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  XOR2_X1   g646(.A(KEYINPUT120), .B(G120gat), .Z(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n840_), .B2(new_n581_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n606_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT121), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n827_), .B(new_n853_), .C1(new_n852_), .C2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g656(.A(new_n842_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT119), .B(new_n838_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n598_), .A2(G127gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G127gat), .B1(new_n827_), .B2(new_n598_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  INV_X1    g663(.A(new_n862_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n864_), .B(new_n865_), .C1(new_n844_), .C2(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n844_), .B2(new_n652_), .ZN(new_n868_));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n827_), .A2(new_n869_), .A3(new_n610_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1343gat));
  NAND3_X1  g670(.A1(new_n659_), .A2(new_n405_), .A3(new_n395_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n825_), .A2(new_n355_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n457_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n606_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n598_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(new_n883_), .A3(new_n610_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n873_), .A2(new_n651_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT125), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n659_), .A2(new_n356_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n646_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n836_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n458_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT22), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n888_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n235_), .B1(new_n893_), .B2(new_n888_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1348gat));
  OR2_X1    g697(.A1(new_n825_), .A2(new_n395_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n659_), .B(new_n356_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n899_), .A2(new_n900_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(G176gat), .A3(new_n606_), .A4(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n904_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n891_), .B2(new_n606_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n892_), .A2(new_n243_), .A3(new_n666_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n901_), .A2(new_n598_), .A3(new_n902_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n222_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n892_), .B2(new_n652_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n891_), .A2(new_n242_), .A3(new_n610_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1351gat));
  NOR2_X1   g713(.A1(new_n825_), .A2(new_n355_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n659_), .A2(new_n411_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n457_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n581_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n207_), .ZN(G1353gat));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n598_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AND2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n923_), .B2(new_n924_), .ZN(G1354gat));
  OAI21_X1  g726(.A(G218gat), .B1(new_n917_), .B2(new_n652_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n623_), .A2(G218gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n917_), .B2(new_n929_), .ZN(G1355gat));
endmodule


