//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  XOR2_X1   g000(.A(G120gat), .B(G148gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G176gat), .B(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT70), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT8), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n211_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n214_), .A3(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n228_));
  INV_X1    g027(.A(G85gat), .ZN(new_n229_));
  INV_X1    g028(.A(G92gat), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT9), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n228_), .A3(new_n231_), .A4(new_n214_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G78gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n224_), .A2(new_n232_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT64), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n224_), .A2(new_n232_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  INV_X1    g050(.A(new_n244_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n241_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n232_), .B(KEYINPUT66), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n224_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT12), .A3(new_n247_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n245_), .A2(new_n250_), .A3(new_n253_), .A4(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n248_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n244_), .B1(new_n258_), .B2(new_n242_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT71), .B(new_n207_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n207_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n260_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n262_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n263_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT13), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n264_), .B(KEYINPUT13), .C1(new_n269_), .C2(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277_));
  INV_X1    g076(.A(G1gat), .ZN(new_n278_));
  INV_X1    g077(.A(G8gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT14), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G43gat), .B(G50gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G29gat), .B(G36gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n283_), .B(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n283_), .A2(new_n289_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n289_), .B(KEYINPUT15), .Z(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  MUX2_X1   g093(.A(new_n290_), .B(new_n293_), .S(new_n294_), .Z(new_n295_));
  XNOR2_X1  g094(.A(G113gat), .B(G141gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT78), .ZN(new_n297_));
  XOR2_X1   g096(.A(G169gat), .B(G197gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT77), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n295_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n276_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT0), .ZN(new_n306_));
  INV_X1    g105(.A(G57gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G85gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(KEYINPUT1), .B2(new_n310_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318_));
  OAI22_X1  g117(.A1(new_n318_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT3), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT2), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n318_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n316_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .A4(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n310_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(new_n311_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n328_), .A2(KEYINPUT86), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT86), .B1(new_n328_), .B2(new_n330_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n317_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n317_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n333_), .A2(new_n343_), .A3(new_n337_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n309_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT96), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n338_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n342_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n346_), .B(new_n309_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT96), .B1(new_n354_), .B2(new_n347_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT22), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G169gat), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n362_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT23), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(G183gat), .A3(G190gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT81), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n370_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n369_), .A2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n370_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT80), .B1(new_n370_), .B2(KEYINPUT23), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n373_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n363_), .A2(new_n367_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n360_), .A2(new_n383_), .A3(KEYINPUT24), .A4(new_n361_), .ZN(new_n384_));
  INV_X1    g183(.A(G183gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT25), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT26), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G190gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n386_), .A2(new_n388_), .A3(new_n390_), .A4(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n383_), .A2(KEYINPUT24), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n382_), .A2(new_n384_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G15gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT82), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n357_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n409_), .A3(new_n357_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n336_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n337_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT21), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT21), .ZN(new_n420_));
  INV_X1    g219(.A(G211gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(G218gat), .ZN(new_n422_));
  INV_X1    g221(.A(G218gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(G211gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n420_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n426_), .A3(KEYINPUT21), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n333_), .B2(KEYINPUT29), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n431_), .B(new_n435_), .C1(new_n333_), .C2(KEYINPUT29), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n417_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n317_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n328_), .A2(new_n330_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n328_), .A2(KEYINPUT86), .A3(new_n330_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n430_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n435_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n432_), .A2(new_n436_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n417_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n439_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G22gat), .B(G50gat), .ZN(new_n455_));
  OR3_X1    g254(.A1(new_n333_), .A2(KEYINPUT29), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(new_n446_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n439_), .A2(KEYINPUT89), .A3(new_n451_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n463_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n416_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n477_));
  AND2_X1   g276(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n478_));
  NOR2_X1   g277(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n383_), .B(new_n358_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n393_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT91), .ZN(new_n482_));
  INV_X1    g281(.A(new_n479_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G169gat), .A2(G176gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n486_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n393_), .A2(new_n480_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n382_), .A2(new_n377_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n369_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n477_), .B1(new_n493_), .B2(new_n430_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n431_), .A2(new_n379_), .A3(new_n395_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n476_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n477_), .B1(new_n396_), .B2(new_n430_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n490_), .A2(new_n431_), .A3(new_n492_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n497_), .A2(new_n476_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n496_), .A2(new_n499_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n362_), .A2(new_n368_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n393_), .A2(new_n480_), .A3(new_n488_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n488_), .B1(new_n393_), .B2(new_n480_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n511_), .B2(new_n487_), .ZN(new_n512_));
  OAI211_X1 g311(.A(KEYINPUT20), .B(new_n495_), .C1(new_n512_), .C2(new_n431_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n475_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n497_), .A2(new_n476_), .A3(new_n498_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n504_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n473_), .B1(new_n506_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n505_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n431_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n521_));
  AND4_X1   g320(.A1(new_n379_), .A2(new_n395_), .A3(new_n429_), .A4(new_n428_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n477_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n515_), .B(new_n504_), .C1(new_n523_), .C2(new_n476_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT98), .A3(new_n473_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n493_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT95), .B1(new_n490_), .B2(new_n492_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n431_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n476_), .B1(new_n531_), .B2(new_n497_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n513_), .A2(new_n475_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n505_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT27), .A3(new_n524_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n472_), .B1(new_n527_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT98), .B1(new_n525_), .B2(new_n473_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n473_), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n518_), .B(new_n538_), .C1(new_n520_), .C2(new_n524_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n472_), .B(new_n535_), .C1(new_n537_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n356_), .B(new_n471_), .C1(new_n536_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT100), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n535_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT99), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT100), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n356_), .A4(new_n471_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n416_), .B(KEYINPUT83), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n466_), .A2(new_n355_), .A3(new_n353_), .A4(new_n470_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(new_n544_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n525_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n309_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n338_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT94), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n354_), .A2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n352_), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n552_), .B(new_n559_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n504_), .A2(KEYINPUT32), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n533_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n497_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n493_), .B(new_n528_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(new_n431_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n569_), .B2(new_n476_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n565_), .B1(new_n570_), .B2(new_n564_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n347_), .B2(new_n354_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n563_), .A2(new_n572_), .B1(new_n470_), .B2(new_n466_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n549_), .B1(new_n551_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n543_), .A2(new_n548_), .A3(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n224_), .A2(new_n232_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT73), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n255_), .B2(new_n292_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(new_n581_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT74), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT75), .B1(new_n590_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n588_), .A2(new_n598_), .A3(new_n595_), .A4(new_n589_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n593_), .B(KEYINPUT36), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n590_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n588_), .A2(KEYINPUT76), .A3(new_n589_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(new_n602_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT76), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n590_), .A2(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n606_), .A2(new_n608_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n609_), .B2(KEYINPUT37), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n283_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n247_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  XOR2_X1   g414(.A(G127gat), .B(G155gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT16), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n614_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(KEYINPUT17), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n304_), .A2(new_n575_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n356_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n278_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT101), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n548_), .A2(new_n574_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n413_), .A2(new_n415_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n465_), .A2(new_n464_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT89), .B1(new_n439_), .B2(new_n451_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n470_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n545_), .B2(new_n540_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n547_), .B1(new_n640_), .B2(new_n356_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n633_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n609_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n276_), .A2(new_n623_), .A3(new_n303_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT102), .Z(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n627_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n631_), .B(new_n632_), .C1(new_n278_), .C2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n546_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n609_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n644_), .A2(new_n649_), .A3(new_n650_), .A4(new_n575_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G8gat), .B1(new_n651_), .B2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT39), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n653_), .A2(new_n654_), .A3(KEYINPUT39), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT104), .B(KEYINPUT39), .C1(new_n653_), .C2(new_n654_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n626_), .A2(new_n279_), .A3(new_n649_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n660_), .A2(KEYINPUT40), .A3(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  INV_X1    g465(.A(new_n549_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n400_), .B1(new_n646_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n626_), .A2(new_n400_), .A3(new_n667_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n637_), .A2(new_n638_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT105), .Z(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n646_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n626_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  INV_X1    g481(.A(new_n623_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n650_), .B2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n609_), .A2(KEYINPUT107), .A3(new_n623_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n304_), .A2(new_n686_), .A3(new_n575_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n627_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n610_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n642_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n575_), .A2(new_n692_), .A3(new_n610_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n274_), .A2(new_n623_), .A3(new_n302_), .A4(new_n275_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT106), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(G29gat), .A3(new_n627_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n696_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n689_), .B1(new_n698_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n649_), .A2(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n649_), .A2(KEYINPUT108), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n688_), .B2(new_n708_), .ZN(new_n709_));
  NOR4_X1   g508(.A1(new_n687_), .A2(new_n707_), .A3(KEYINPUT45), .A4(G36gat), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n709_), .A2(new_n710_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n701_), .A2(new_n649_), .A3(new_n697_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(G36gat), .ZN(new_n713_));
  AND2_X1   g512(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n701_), .A2(G43gat), .A3(new_n634_), .A4(new_n697_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n687_), .A2(new_n549_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(G43gat), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g518(.A(G50gat), .B1(new_n688_), .B2(new_n676_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n697_), .A2(G50gat), .A3(new_n675_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n701_), .ZN(G1331gat));
  AOI211_X1 g521(.A(new_n623_), .B(new_n302_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n643_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n643_), .A2(new_n723_), .A3(KEYINPUT112), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G57gat), .A3(new_n627_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n624_), .A2(new_n276_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT110), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n303_), .C1(new_n633_), .C2(new_n641_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n303_), .B1(new_n633_), .B2(new_n641_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n627_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n730_), .A2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n728_), .B2(new_n706_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(new_n740_), .A3(new_n706_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n728_), .B2(new_n667_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n737_), .A2(new_n745_), .A3(new_n667_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n737_), .A2(new_n750_), .A3(new_n676_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n726_), .A2(new_n676_), .A3(new_n727_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G78gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G78gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1335gat));
  NAND3_X1  g557(.A1(new_n276_), .A2(new_n623_), .A3(new_n303_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n356_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n276_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n685_), .B2(new_n684_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n734_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n733_), .B1(new_n575_), .B2(new_n303_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT115), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n736_), .A2(new_n734_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n764_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n627_), .A2(new_n229_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n762_), .B1(new_n773_), .B2(new_n774_), .ZN(G1336gat));
  OAI21_X1  g574(.A(G92gat), .B1(new_n761_), .B2(new_n707_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n649_), .A2(new_n230_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(G1337gat));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n634_), .A2(new_n225_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n769_), .B2(new_n764_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n686_), .A2(new_n276_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT115), .B(new_n783_), .C1(new_n736_), .C2(new_n734_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n760_), .A2(new_n667_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G99gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n785_), .A2(new_n786_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n780_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n791_));
  INV_X1    g590(.A(G99gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n760_), .B2(new_n667_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT51), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n772_), .B2(new_n781_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n786_), .B1(new_n796_), .B2(new_n789_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n779_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n785_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n800_), .A2(KEYINPUT118), .A3(new_n790_), .A4(new_n794_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n772_), .A2(new_n226_), .A3(new_n675_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n760_), .A2(new_n675_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G106gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT52), .B(new_n226_), .C1(new_n760_), .C2(new_n675_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g608(.A(new_n302_), .B1(new_n207_), .B2(new_n260_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n250_), .A2(new_n256_), .A3(new_n241_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n244_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT119), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n257_), .B(KEYINPUT55), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n265_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT120), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n816_), .B2(KEYINPUT56), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n815_), .B2(KEYINPUT120), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n295_), .A2(new_n300_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n293_), .A2(G229gat), .A3(G233gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n290_), .A2(new_n294_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n300_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n272_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT57), .B(new_n650_), .C1(new_n820_), .C2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n817_), .A2(new_n819_), .B1(new_n272_), .B2(new_n826_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n609_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n815_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  INV_X1    g633(.A(new_n815_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n818_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n833_), .B(new_n836_), .C1(KEYINPUT56), .C2(new_n815_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n825_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT58), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n838_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n610_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n683_), .B1(new_n832_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n763_), .A2(new_n303_), .A3(new_n624_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT54), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n627_), .B(new_n640_), .C1(new_n843_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n610_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n831_), .B(new_n828_), .C1(new_n850_), .C2(new_n839_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n623_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n845_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n853_), .A2(KEYINPUT59), .A3(new_n627_), .A4(new_n640_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n303_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n302_), .A2(new_n856_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n855_), .A2(new_n856_), .B1(new_n847_), .B2(new_n857_), .ZN(G1340gat));
  AOI21_X1  g657(.A(new_n763_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT122), .B(G120gat), .Z(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n763_), .A2(KEYINPUT60), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(KEYINPUT60), .B2(new_n861_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n859_), .A2(new_n860_), .B1(new_n847_), .B2(new_n863_), .ZN(G1341gat));
  AOI21_X1  g663(.A(new_n623_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n865_));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n683_), .A2(new_n866_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n865_), .A2(new_n866_), .B1(new_n847_), .B2(new_n867_), .ZN(G1342gat));
  NAND2_X1  g667(.A1(new_n849_), .A2(new_n854_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n610_), .A2(G134gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT123), .Z(new_n871_));
  OR2_X1    g670(.A1(new_n847_), .A2(new_n650_), .ZN(new_n872_));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n869_), .A2(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1343gat));
  NOR4_X1   g673(.A1(new_n706_), .A2(new_n638_), .A3(new_n637_), .A4(new_n667_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n853_), .A2(new_n627_), .A3(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n303_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT124), .B(G141gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1344gat));
  OR3_X1    g678(.A1(new_n876_), .A2(G148gat), .A3(new_n763_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G148gat), .B1(new_n876_), .B2(new_n763_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1345gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n876_), .A2(new_n623_), .A3(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n876_), .B2(new_n623_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n876_), .B2(new_n690_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n650_), .A2(G162gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n876_), .B2(new_n889_), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n707_), .A2(new_n627_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n667_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n676_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n853_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n302_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT125), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n853_), .A2(new_n302_), .A3(new_n893_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n894_), .B2(new_n276_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n843_), .A2(new_n846_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n675_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n892_), .A2(new_n367_), .A3(new_n763_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  NAND4_X1  g706(.A1(new_n905_), .A2(new_n667_), .A3(new_n683_), .A4(new_n891_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n623_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n908_), .A2(new_n385_), .B1(new_n894_), .B2(new_n909_), .ZN(G1350gat));
  NAND4_X1  g709(.A1(new_n894_), .A2(new_n609_), .A3(new_n390_), .A4(new_n392_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n894_), .A2(new_n610_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n389_), .ZN(G1351gat));
  NAND3_X1  g712(.A1(new_n891_), .A2(new_n675_), .A3(new_n549_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n904_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n302_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  XOR2_X1   g716(.A(KEYINPUT126), .B(G204gat), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n915_), .B2(new_n276_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n915_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n763_), .ZN(new_n921_));
  INV_X1    g720(.A(G204gat), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(KEYINPUT126), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n921_), .B2(new_n923_), .ZN(G1353gat));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n683_), .B1(new_n925_), .B2(new_n421_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT127), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n915_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n925_), .A2(new_n421_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n920_), .B2(new_n690_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n915_), .A2(new_n423_), .A3(new_n609_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


