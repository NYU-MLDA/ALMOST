//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT66), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT67), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n214_), .A2(new_n216_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G29gat), .B(G36gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT68), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n232_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT7), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n233_), .A2(new_n235_), .A3(new_n238_), .A4(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n209_), .A2(new_n212_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(KEYINPUT70), .A3(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n223_), .A2(new_n217_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n230_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n214_), .B2(new_n243_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n226_), .B(new_n229_), .C1(new_n251_), .C2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT77), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n258_), .A2(new_n260_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT80), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n255_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n226_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n229_), .B(KEYINPUT15), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT75), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n247_), .A2(new_n246_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT70), .B1(new_n241_), .B2(new_n242_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n250_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n246_), .A2(KEYINPUT67), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n213_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n274_), .A3(new_n243_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n271_), .A2(KEYINPUT8), .B1(new_n275_), .B2(new_n252_), .ZN(new_n276_));
  AND4_X1   g075(.A1(new_n216_), .A2(new_n272_), .A3(new_n274_), .A4(new_n225_), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT75), .B(new_n267_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n265_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT76), .B1(new_n279_), .B2(new_n268_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n255_), .A2(new_n262_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n271_), .A2(KEYINPUT8), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n252_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n277_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n267_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n283_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n278_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n263_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n280_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n299_));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G134gat), .B(G162gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n294_), .B1(new_n291_), .B2(new_n263_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT36), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n303_), .A2(new_n305_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n298_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n298_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n202_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n298_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n298_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT37), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT82), .B(G15gat), .ZN(new_n317_));
  INV_X1    g116(.A(G22gat), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT83), .B(G1gat), .ZN(new_n320_));
  INV_X1    g119(.A(G8gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT14), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n318_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G8gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G57gat), .B(G64gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT11), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G71gat), .B(G78gat), .Z(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(KEYINPUT11), .B2(new_n332_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n331_), .B(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G183gat), .B(G211gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G155gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n344_), .A2(KEYINPUT17), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(KEYINPUT17), .B2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n339_), .A2(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT85), .B1(new_n339_), .B2(new_n345_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n347_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n316_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT94), .B(G204gat), .ZN(new_n354_));
  INV_X1    g153(.A(G197gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G204gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n356_), .B(KEYINPUT21), .C1(new_n355_), .C2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(G197gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(G197gat), .B2(new_n357_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n358_), .B(new_n359_), .C1(new_n361_), .C2(KEYINPUT21), .ZN(new_n362_));
  INV_X1    g161(.A(new_n359_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(KEYINPUT21), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  OR2_X1    g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT3), .Z(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT2), .Z(new_n371_));
  OAI211_X1 g170(.A(new_n366_), .B(new_n367_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n367_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n373_), .B(new_n370_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n365_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n382_), .A2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n379_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G78gat), .B(G106gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n390_), .A2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n387_), .A2(new_n394_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT0), .B(G57gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT91), .ZN(new_n406_));
  XOR2_X1   g205(.A(G113gat), .B(G120gat), .Z(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n407_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT92), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n406_), .A2(KEYINPUT92), .A3(new_n407_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n378_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(KEYINPUT96), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT96), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n409_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(new_n378_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT4), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n412_), .A2(KEYINPUT4), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n404_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(KEYINPUT96), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n404_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n403_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n419_), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n427_), .B(new_n402_), .C1(new_n428_), .C2(new_n404_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G183gat), .ZN(new_n431_));
  INV_X1    g230(.A(G190gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT23), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT88), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G183gat), .A3(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(G183gat), .B2(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G169gat), .A2(G176gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G169gat), .ZN(new_n440_));
  INV_X1    g239(.A(G176gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n436_), .A2(KEYINPUT90), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(KEYINPUT90), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n433_), .A3(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT24), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT95), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n447_), .A2(new_n439_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT25), .B(G183gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT26), .B(G190gat), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n452_), .A2(KEYINPUT24), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(KEYINPUT95), .A3(new_n448_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n443_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n365_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n442_), .A2(new_n439_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT89), .Z(new_n461_));
  OAI21_X1  g260(.A(new_n446_), .B1(G183gat), .B2(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n437_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n459_), .B(KEYINPUT20), .C1(new_n465_), .C2(new_n365_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G226gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT19), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n443_), .A2(new_n362_), .A3(new_n364_), .A4(new_n457_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT20), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n465_), .B2(new_n365_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n222_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT18), .B(G64gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OR3_X1    g281(.A1(new_n475_), .A2(KEYINPUT98), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n468_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n472_), .A2(KEYINPUT99), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT99), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n471_), .A2(new_n486_), .B1(new_n465_), .B2(new_n365_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n484_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n466_), .A2(new_n468_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n482_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT98), .B1(new_n475_), .B2(new_n482_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n430_), .A2(new_n483_), .A3(new_n490_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n429_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n421_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(KEYINPUT33), .A3(new_n402_), .A4(new_n427_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n469_), .A2(new_n480_), .A3(new_n474_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n480_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n403_), .B1(new_n423_), .B2(new_n404_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT97), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT97), .B(new_n403_), .C1(new_n423_), .C2(new_n404_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n503_), .B(new_n504_), .C1(new_n424_), .C2(new_n428_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n494_), .A2(new_n496_), .A3(new_n500_), .A4(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n398_), .B1(new_n492_), .B2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n410_), .A2(new_n411_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT31), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n508_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n465_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G99gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G43gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT30), .B(G15gat), .Z(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n397_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n526_), .A2(new_n522_), .A3(new_n521_), .A4(new_n395_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n426_), .A2(new_n429_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT27), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n479_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT27), .A3(new_n497_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n529_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n507_), .A2(new_n524_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n338_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n226_), .B(new_n338_), .C1(new_n251_), .C2(new_n254_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(KEYINPUT12), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n266_), .A2(new_n540_), .A3(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT64), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n537_), .A2(new_n538_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT5), .B(G176gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G204gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n550_), .B(KEYINPUT72), .ZN(new_n559_));
  INV_X1    g358(.A(new_n557_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n546_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n561_), .A3(KEYINPUT13), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n329_), .A2(new_n229_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n287_), .B2(new_n329_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n568_), .A2(KEYINPUT86), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n329_), .B(new_n229_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT86), .B1(new_n568_), .B2(new_n570_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT87), .B(G113gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .A4(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n566_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n535_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n353_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(new_n430_), .A3(new_n320_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT38), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT100), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(KEYINPUT38), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n313_), .A2(new_n314_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n352_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n585_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n529_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n596_), .ZN(G1324gat));
  AND2_X1   g396(.A1(new_n533_), .A2(new_n531_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G8gat), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT39), .ZN(new_n600_));
  INV_X1    g399(.A(new_n598_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n587_), .A2(new_n321_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g403(.A(G15gat), .B1(new_n595_), .B2(new_n524_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n586_), .A2(G15gat), .A3(new_n524_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT101), .Z(G1326gat));
  XOR2_X1   g408(.A(new_n398_), .B(KEYINPUT102), .Z(new_n610_));
  OAI21_X1  g409(.A(G22gat), .B1(new_n595_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT42), .ZN(new_n612_));
  INV_X1    g411(.A(new_n610_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n587_), .A2(new_n318_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1327gat));
  INV_X1    g414(.A(new_n352_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n592_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n585_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n585_), .A2(new_n617_), .A3(KEYINPUT105), .ZN(new_n621_));
  INV_X1    g420(.A(G29gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n430_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT106), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n310_), .A2(new_n315_), .B1(new_n535_), .B2(KEYINPUT103), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n535_), .A2(KEYINPUT103), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n535_), .A2(KEYINPUT43), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n316_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n316_), .B2(new_n632_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n630_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n584_), .A2(new_n616_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n626_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n634_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n316_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n628_), .A2(new_n629_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n639_), .B(new_n640_), .C1(new_n641_), .C2(new_n627_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n636_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n638_), .A2(new_n643_), .A3(new_n430_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n625_), .B1(new_n644_), .B2(new_n622_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT107), .B(new_n625_), .C1(new_n644_), .C2(new_n622_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n620_), .A2(new_n650_), .A3(new_n601_), .A4(new_n621_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n638_), .A2(new_n643_), .A3(new_n601_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(G36gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT108), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT108), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  NAND4_X1  g460(.A1(new_n638_), .A2(new_n643_), .A3(G43gat), .A4(new_n523_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT109), .B(G43gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n620_), .A2(new_n621_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n524_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g466(.A1(new_n638_), .A2(new_n643_), .A3(new_n398_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT110), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT110), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(G50gat), .A3(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n610_), .A2(G50gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n664_), .B2(new_n672_), .ZN(G1331gat));
  NOR2_X1   g472(.A1(new_n566_), .A2(new_n583_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n535_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n353_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT111), .ZN(new_n678_));
  AOI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n430_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n594_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n529_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(G57gat), .B2(new_n681_), .ZN(G1332gat));
  INV_X1    g481(.A(G64gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(new_n683_), .A3(new_n601_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G64gat), .B1(new_n680_), .B2(new_n598_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT48), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1333gat));
  INV_X1    g486(.A(G71gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n678_), .A2(new_n688_), .A3(new_n523_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G71gat), .B1(new_n680_), .B2(new_n524_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT49), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1334gat));
  INV_X1    g491(.A(G78gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n693_), .A3(new_n613_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G78gat), .B1(new_n680_), .B2(new_n610_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT50), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1335gat));
  NOR3_X1   g496(.A1(new_n635_), .A2(new_n616_), .A3(new_n675_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G85gat), .A3(new_n430_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n676_), .A2(new_n617_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n221_), .B1(new_n700_), .B2(new_n529_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1336gat));
  NAND3_X1  g501(.A1(new_n698_), .A2(G92gat), .A3(new_n601_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n222_), .B1(new_n700_), .B2(new_n598_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1337gat));
  NOR3_X1   g504(.A1(new_n700_), .A2(new_n215_), .A3(new_n524_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(new_n523_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G99gat), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT51), .Z(G1338gat));
  NOR2_X1   g508(.A1(new_n675_), .A2(new_n616_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n642_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n398_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G106gat), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(KEYINPUT114), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(KEYINPUT114), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n713_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n700_), .A2(G106gat), .A3(new_n712_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(new_n721_));
  OAI211_X1 g520(.A(G106gat), .B(new_n716_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT53), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n719_), .A2(new_n725_), .A3(new_n721_), .A4(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(new_n583_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n564_), .A2(new_n616_), .A3(new_n728_), .A4(new_n565_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT115), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n572_), .A2(new_n569_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n580_), .C1(new_n569_), .C2(new_n568_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n582_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT55), .B1(new_n542_), .B2(new_n545_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n546_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n542_), .A2(KEYINPUT55), .A3(new_n545_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n542_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n545_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n557_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n561_), .B(new_n737_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT58), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n744_), .A2(new_n557_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT58), .A3(new_n561_), .A4(new_n737_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n308_), .A2(new_n309_), .A3(new_n202_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT37), .B1(new_n313_), .B2(new_n314_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n749_), .B(new_n755_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n561_), .A2(new_n583_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n553_), .A2(new_n557_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n560_), .B1(new_n559_), .B2(new_n546_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n737_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n562_), .A2(KEYINPUT118), .A3(new_n737_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n761_), .A2(new_n768_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT118), .B1(new_n562_), .B2(new_n737_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n765_), .B(new_n736_), .C1(new_n558_), .C2(new_n561_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n760_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n592_), .A3(KEYINPUT57), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n758_), .A2(new_n759_), .A3(new_n771_), .A4(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n352_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n777_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT57), .B1(new_n777_), .B2(new_n592_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n759_), .B1(new_n783_), .B2(new_n758_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n733_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n601_), .A2(new_n529_), .A3(new_n525_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n583_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n749_), .A2(new_n755_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n315_), .B2(new_n310_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n771_), .A2(new_n778_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n352_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT120), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n352_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n733_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n786_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n790_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n728_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n789_), .B1(new_n802_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n801_), .B2(new_n566_), .ZN(new_n804_));
  INV_X1    g603(.A(G120gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n788_), .B(new_n806_), .C1(KEYINPUT60), .C2(new_n805_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n788_), .B2(new_n616_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n790_), .A2(G127gat), .A3(new_n800_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n616_), .ZN(G1342gat));
  AOI21_X1  g610(.A(G134gat), .B1(new_n788_), .B2(new_n593_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n801_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n316_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT121), .B(G134gat), .Z(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT122), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n813_), .B2(new_n817_), .ZN(G1343gat));
  AND3_X1   g617(.A1(new_n785_), .A2(new_n524_), .A3(new_n398_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n601_), .A2(new_n529_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n583_), .A3(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g621(.A(new_n566_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n823_), .A3(new_n820_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g624(.A1(new_n819_), .A2(new_n616_), .A3(new_n820_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  AND4_X1   g627(.A1(G162gat), .A2(new_n819_), .A3(new_n316_), .A4(new_n820_), .ZN(new_n829_));
  INV_X1    g628(.A(G162gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(new_n593_), .A3(new_n820_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(G1347gat));
  NOR2_X1   g631(.A1(new_n598_), .A2(new_n430_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n523_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT123), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n798_), .A2(new_n610_), .A3(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G169gat), .B1(new_n836_), .B2(new_n728_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n798_), .A2(new_n610_), .A3(new_n835_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n583_), .A3(new_n440_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(G1348gat));
  AND3_X1   g642(.A1(new_n835_), .A2(G176gat), .A3(new_n823_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n785_), .A2(KEYINPUT124), .A3(new_n712_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT124), .B1(new_n785_), .B2(new_n712_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT125), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n441_), .B1(new_n836_), .B2(new_n566_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n844_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n848_), .A2(new_n849_), .A3(new_n851_), .ZN(G1349gat));
  NAND2_X1  g651(.A1(new_n785_), .A2(new_n712_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n785_), .A2(KEYINPUT124), .A3(new_n712_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n352_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G183gat), .B1(new_n857_), .B2(new_n835_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  INV_X1    g658(.A(new_n453_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n840_), .A2(new_n859_), .A3(new_n616_), .A4(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n798_), .A2(new_n860_), .A3(new_n610_), .A4(new_n835_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT126), .B1(new_n862_), .B2(new_n352_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n858_), .A2(new_n864_), .ZN(G1350gat));
  AOI21_X1  g664(.A(new_n432_), .B1(new_n840_), .B2(new_n316_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n798_), .A2(new_n454_), .A3(new_n610_), .A4(new_n835_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n592_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT127), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G190gat), .B1(new_n836_), .B2(new_n814_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT127), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n870_), .B(new_n871_), .C1(new_n592_), .C2(new_n867_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(G1351gat));
  NAND3_X1  g672(.A1(new_n819_), .A2(new_n583_), .A3(new_n833_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g674(.A1(new_n819_), .A2(new_n833_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n823_), .A3(new_n354_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n819_), .A2(new_n833_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G204gat), .B1(new_n878_), .B2(new_n566_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1353gat));
  NAND3_X1  g679(.A1(new_n819_), .A2(new_n616_), .A3(new_n833_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT63), .B(G211gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n881_), .B2(new_n884_), .ZN(G1354gat));
  AOI21_X1  g684(.A(G218gat), .B1(new_n876_), .B2(new_n593_), .ZN(new_n886_));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n878_), .A2(new_n887_), .A3(new_n814_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1355gat));
endmodule


