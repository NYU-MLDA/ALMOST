//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  OR3_X1    g007(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n203_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT22), .B(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n205_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n205_), .B1(new_n216_), .B2(KEYINPUT22), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G169gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(KEYINPUT81), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT81), .B1(new_n217_), .B2(new_n219_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G227gat), .A2(G233gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n225_), .B(KEYINPUT82), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G99gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G134gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G127gat), .ZN(new_n234_));
  INV_X1    g033(.A(G127gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G134gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT83), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n232_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(KEYINPUT83), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n231_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT31), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G15gat), .B(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n230_), .B(new_n249_), .Z(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  XOR2_X1   g051(.A(G211gat), .B(G218gat), .Z(new_n253_));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254_));
  INV_X1    g053(.A(G204gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(G197gat), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n253_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT90), .B1(new_n255_), .B2(G197gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n257_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n255_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT21), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n253_), .A2(KEYINPUT21), .ZN(new_n268_));
  INV_X1    g067(.A(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n224_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n211_), .A2(KEYINPUT93), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n211_), .A2(KEYINPUT93), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n212_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n207_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n215_), .B2(new_n205_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n275_), .A2(new_n210_), .B1(new_n221_), .B2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n262_), .A2(new_n266_), .B1(new_n269_), .B2(new_n268_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n252_), .B1(new_n272_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G8gat), .B(G36gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n224_), .A2(new_n271_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n252_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n279_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n286_), .A2(KEYINPUT20), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT27), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(KEYINPUT20), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT97), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n292_), .A2(KEYINPUT97), .B1(new_n224_), .B2(new_n271_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n272_), .A2(new_n280_), .A3(new_n252_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n285_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n291_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n281_), .A2(KEYINPUT94), .A3(new_n289_), .A4(new_n285_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n281_), .A2(new_n289_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n285_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n290_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT100), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n290_), .A2(new_n304_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n301_), .C1(new_n285_), .C2(new_n302_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT100), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n300_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n299_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT84), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n317_), .A2(new_n314_), .A3(new_n315_), .A4(KEYINPUT84), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n319_), .A2(new_n320_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n316_), .A2(new_n321_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(KEYINPUT1), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G155gat), .A3(G162gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n333_), .A3(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n246_), .A2(new_n336_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n325_), .A2(new_n328_), .B1(new_n334_), .B2(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT4), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n246_), .A2(new_n336_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n313_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  INV_X1    g143(.A(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n313_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n343_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n348_), .B1(new_n343_), .B2(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT98), .B(new_n348_), .C1(new_n343_), .C2(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G106gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n336_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT88), .B1(new_n362_), .B2(new_n358_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n338_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(new_n279_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(G78gat), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n359_), .A2(new_n360_), .B1(G228gat), .B2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n357_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(G78gat), .A3(new_n368_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n371_), .B1(new_n370_), .B2(new_n367_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(G106gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(KEYINPUT87), .A3(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G22gat), .B(G50gat), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n338_), .A2(new_n365_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT86), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n375_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n357_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n378_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n376_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n383_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n377_), .A2(new_n378_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n386_), .B2(new_n376_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n312_), .A2(new_n356_), .A3(new_n389_), .A4(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT101), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n389_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n353_), .A2(KEYINPUT33), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n348_), .C1(new_n343_), .C2(new_n350_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n340_), .A2(new_n313_), .A3(new_n342_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n403_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n337_), .A2(new_n339_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n348_), .B1(new_n406_), .B2(new_n349_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT96), .B1(new_n409_), .B2(new_n309_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n303_), .A2(new_n305_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n401_), .A4(new_n408_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT32), .B(new_n285_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT32), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n302_), .B1(new_n415_), .B2(new_n298_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n414_), .A2(new_n355_), .A3(new_n354_), .A4(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n397_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT99), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n379_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n383_), .B1(new_n379_), .B2(new_n388_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n423_), .A2(KEYINPUT101), .A3(new_n356_), .A4(new_n312_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT99), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n397_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n396_), .A2(new_n420_), .A3(new_n424_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT102), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n397_), .A2(new_n428_), .A3(new_n312_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n397_), .B2(new_n312_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n250_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n250_), .A2(new_n427_), .B1(new_n431_), .B2(new_n356_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT36), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G232gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT72), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT64), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT9), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G92gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT64), .B1(new_n345_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n441_), .B(new_n444_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n357_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n357_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT15), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n439_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n448_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n450_), .A2(new_n452_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n458_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n464_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT8), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n473_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n470_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n480_), .A2(KEYINPUT71), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(KEYINPUT71), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n472_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n436_), .A2(new_n437_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G190gat), .B(G218gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT73), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G134gat), .B(G162gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  OAI221_X1 g288(.A(new_n472_), .B1(new_n437_), .B2(new_n436_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n490_));
  AND4_X1   g289(.A1(new_n433_), .A2(new_n485_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n489_), .B(new_n433_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n432_), .A2(KEYINPUT104), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT104), .B1(new_n432_), .B2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G57gat), .ZN(new_n505_));
  INV_X1    g304(.A(G57gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G64gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n502_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n457_), .B(new_n511_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n479_), .B2(new_n511_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n499_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT12), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(KEYINPUT12), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n479_), .B2(new_n511_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n511_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n467_), .A2(new_n523_), .A3(new_n520_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n519_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n498_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G120gat), .B(G148gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n516_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n526_), .B2(new_n516_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT13), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n470_), .B(KEYINPUT76), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540_));
  INV_X1    g339(.A(G1gat), .ZN(new_n541_));
  INV_X1    g340(.A(G8gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G1gat), .B(G8gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT77), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n471_), .A2(new_n546_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n539_), .A2(new_n546_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n556_), .B2(new_n550_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT79), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  OAI221_X1 g361(.A(new_n552_), .B1(KEYINPUT79), .B2(new_n560_), .C1(new_n556_), .C2(new_n550_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n538_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT103), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n546_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n523_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT16), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n569_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n569_), .A2(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n569_), .A2(KEYINPUT75), .A3(new_n575_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n566_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n497_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n356_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n427_), .A2(new_n250_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n431_), .A2(new_n356_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n538_), .B(KEYINPUT68), .ZN(new_n590_));
  OR2_X1    g389(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n591_));
  NAND2_X1  g390(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n591_), .B(new_n592_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n493_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n485_), .A2(new_n433_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n594_), .A2(KEYINPUT74), .A3(KEYINPUT37), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n582_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n590_), .A2(new_n564_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n589_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n356_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n541_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n586_), .A2(new_n604_), .ZN(G1324gat));
  XNOR2_X1  g404(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT106), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n312_), .B(new_n583_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n542_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT106), .B(G8gat), .C1(new_n585_), .C2(new_n312_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT39), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n608_), .B(new_n613_), .C1(new_n609_), .C2(new_n542_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n312_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n542_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT105), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n607_), .B1(new_n612_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT39), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(new_n614_), .A3(new_n617_), .A4(new_n606_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1325gat));
  INV_X1    g421(.A(new_n601_), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n623_), .A2(G15gat), .A3(new_n250_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n250_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n497_), .A2(new_n625_), .A3(new_n584_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(new_n626_), .B2(G15gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(G1326gat));
  OR3_X1    g428(.A1(new_n623_), .A2(G22gat), .A3(new_n397_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n497_), .A2(new_n423_), .A3(new_n584_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT42), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G22gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G22gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(new_n494_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n432_), .A2(new_n636_), .A3(new_n582_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n565_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n602_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n597_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n589_), .B2(new_n597_), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n598_), .B(new_n642_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n582_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n566_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT109), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n646_), .C2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n602_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n639_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NOR2_X1   g454(.A1(new_n312_), .A2(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n637_), .A2(new_n565_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT110), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n637_), .A2(new_n659_), .A3(new_n565_), .A4(new_n656_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(KEYINPUT45), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT45), .B1(new_n658_), .B2(new_n660_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n312_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n664_));
  INV_X1    g463(.A(G36gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n663_), .B(KEYINPUT46), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1329gat));
  AOI21_X1  g469(.A(G43gat), .B1(new_n638_), .B2(new_n625_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n625_), .A2(G43gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n653_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1330gat));
  INV_X1    g474(.A(G50gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n638_), .A2(new_n676_), .A3(new_n423_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n653_), .A2(KEYINPUT111), .A3(new_n423_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G50gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT111), .B1(new_n653_), .B2(new_n423_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n562_), .A2(new_n563_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n647_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n590_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n497_), .A2(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n685_), .A2(new_n506_), .A3(new_n356_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n538_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n599_), .A2(new_n682_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n589_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n506_), .B1(new_n689_), .B2(new_n356_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT112), .Z(new_n691_));
  NOR2_X1   g490(.A1(new_n686_), .A2(new_n691_), .ZN(G1332gat));
  INV_X1    g491(.A(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n504_), .A3(new_n615_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  INV_X1    g494(.A(new_n685_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n615_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n697_), .B2(G64gat), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT48), .B(new_n504_), .C1(new_n696_), .C2(new_n615_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1333gat));
  OR3_X1    g499(.A1(new_n689_), .A2(G71gat), .A3(new_n250_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G71gat), .B1(new_n685_), .B2(new_n250_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT49), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT49), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1334gat));
  NAND3_X1  g504(.A1(new_n693_), .A2(new_n371_), .A3(new_n423_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n696_), .A2(new_n423_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G78gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT50), .B(new_n371_), .C1(new_n696_), .C2(new_n423_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n687_), .A2(new_n682_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n647_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n642_), .B1(new_n432_), .B2(new_n598_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n589_), .A2(new_n597_), .A3(new_n643_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n356_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n590_), .A2(new_n564_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n637_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n345_), .A3(new_n602_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n717_), .B2(new_n312_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n445_), .A3(new_n615_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n717_), .B2(new_n250_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n720_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n625_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g529(.A(new_n357_), .B1(new_n716_), .B2(new_n423_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT115), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n713_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n423_), .B(new_n734_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n732_), .A3(G106gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n397_), .B(new_n713_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n739_), .B(KEYINPUT52), .C1(new_n740_), .C2(new_n357_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n735_), .A2(KEYINPUT114), .A3(new_n732_), .A4(G106gat), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n733_), .A2(new_n738_), .A3(new_n741_), .A4(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n720_), .A2(new_n357_), .A3(new_n423_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT113), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n564_), .A2(new_n536_), .A3(new_n582_), .A4(new_n537_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n687_), .A2(new_n754_), .A3(new_n683_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n751_), .B1(new_n756_), .B2(new_n598_), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT54), .B(new_n597_), .C1(new_n753_), .C2(new_n755_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n560_), .B(new_n552_), .C1(new_n556_), .C2(new_n550_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n560_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n549_), .A2(new_n555_), .A3(new_n550_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n550_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n535_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n512_), .A2(new_n518_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n479_), .A2(new_n511_), .A3(new_n521_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n520_), .B1(new_n467_), .B2(new_n523_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n499_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(KEYINPUT55), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n768_), .B(KEYINPUT55), .C1(new_n525_), .C2(new_n498_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n526_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n531_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT55), .B1(new_n525_), .B2(new_n498_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT117), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n780_), .A2(new_n498_), .A3(new_n525_), .A4(new_n775_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n775_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n531_), .B1(new_n787_), .B2(new_n526_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n781_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT118), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n781_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n564_), .A2(new_n533_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n767_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n760_), .B1(new_n794_), .B2(new_n494_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n789_), .B2(KEYINPUT118), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n784_), .A2(new_n785_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n767_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n766_), .A2(new_n533_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n782_), .A2(new_n783_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n789_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n598_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n802_), .B(KEYINPUT58), .C1(new_n803_), .C2(new_n789_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n784_), .A2(new_n791_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n802_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n795_), .A2(new_n801_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n759_), .B1(new_n813_), .B2(new_n647_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n431_), .A2(new_n602_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n682_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n759_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n647_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n813_), .B2(new_n647_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n431_), .A2(KEYINPUT120), .A3(new_n602_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT59), .B1(new_n814_), .B2(new_n815_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n682_), .A2(G113gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT122), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n817_), .B1(new_n831_), .B2(new_n833_), .ZN(G1340gat));
  AOI21_X1  g633(.A(new_n494_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n812_), .B1(new_n835_), .B2(KEYINPUT57), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n794_), .A2(new_n760_), .A3(new_n494_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n647_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n647_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n759_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n590_), .B(new_n829_), .C1(new_n842_), .C2(new_n826_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n828_), .A2(KEYINPUT123), .A3(new_n590_), .A4(new_n829_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(G120gat), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n687_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n816_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT124), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n853_), .A3(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n816_), .B2(new_n582_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n235_), .B1(new_n582_), .B2(KEYINPUT125), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(KEYINPUT125), .B2(new_n235_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n831_), .B2(new_n858_), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n830_), .B2(new_n598_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n816_), .A2(new_n233_), .A3(new_n494_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n814_), .A2(new_n625_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n602_), .A3(new_n423_), .A4(new_n312_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n865_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n682_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g668(.A(new_n590_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g670(.A(new_n582_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  NOR2_X1   g673(.A1(new_n866_), .A2(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G162gat), .B1(new_n875_), .B2(new_n598_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n636_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n312_), .A2(new_n602_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n250_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n842_), .A2(new_n423_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n682_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n204_), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n884_), .B(new_n885_), .C1(KEYINPUT127), .C2(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(new_n215_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n888_), .B(new_n889_), .C1(new_n890_), .C2(new_n884_), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n883_), .B2(new_n538_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n814_), .A2(new_n423_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n881_), .A2(G176gat), .A3(new_n590_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n882_), .A2(new_n647_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G183gat), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n273_), .A2(new_n274_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n582_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n897_), .B1(new_n883_), .B2(new_n900_), .ZN(G1350gat));
  NAND2_X1  g700(.A1(new_n883_), .A2(new_n597_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G190gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n883_), .A2(new_n494_), .A3(new_n212_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n880_), .A2(new_n397_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n863_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n564_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n258_), .ZN(G1352gat));
  INV_X1    g708(.A(new_n907_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n590_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n582_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  OR3_X1    g716(.A1(new_n907_), .A2(G218gat), .A3(new_n636_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G218gat), .B1(new_n907_), .B2(new_n598_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1355gat));
endmodule


