//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_;
  XOR2_X1   g000(.A(G169gat), .B(G197gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT85), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n210_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n211_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(new_n214_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G29gat), .B(G36gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT15), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n216_), .A2(new_n218_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(KEYINPUT83), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT84), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT84), .B1(new_n225_), .B2(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n224_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n226_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n227_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n219_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n231_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n205_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n231_), .A3(new_n224_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n205_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n236_), .A2(new_n227_), .B1(new_n219_), .B2(new_n238_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n242_), .B(new_n243_), .C1(new_n231_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT22), .B(G169gat), .Z(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT87), .B(new_n248_), .C1(new_n249_), .C2(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  OR2_X1    g050(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(G176gat), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n248_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257_));
  INV_X1    g056(.A(G183gat), .ZN(new_n258_));
  INV_X1    g057(.A(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n250_), .A2(new_n256_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT25), .B(G183gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT86), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n259_), .B2(KEYINPUT26), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(KEYINPUT26), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT26), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT86), .A3(G190gat), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n270_), .B(new_n277_), .C1(new_n255_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n264_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G15gat), .B(G43gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT31), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n280_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G71gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n288_), .A2(new_n289_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n285_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n286_), .B(new_n287_), .Z(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G71gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(G227gat), .A3(new_n290_), .A4(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT30), .B(G99gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n293_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n284_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n297_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n283_), .A3(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G22gat), .B(G50gat), .Z(new_n307_));
  INV_X1    g106(.A(G141gat), .ZN(new_n308_));
  INV_X1    g107(.A(G148gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n308_), .B(new_n309_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT88), .B1(new_n321_), .B2(KEYINPUT1), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(G155gat), .A4(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(KEYINPUT1), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .A4(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n310_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n307_), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  INV_X1    g134(.A(new_n307_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n323_), .A2(new_n335_), .A3(new_n331_), .A4(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n334_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT93), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n335_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(G197gat), .ZN(new_n346_));
  INV_X1    g145(.A(G197gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT21), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT92), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n347_), .A3(G204gat), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT92), .B1(new_n345_), .B2(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(new_n346_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n344_), .B(new_n349_), .C1(new_n353_), .C2(KEYINPUT21), .ZN(new_n354_));
  INV_X1    g153(.A(new_n344_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n355_), .A3(KEYINPUT21), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT91), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n343_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n343_), .B2(new_n359_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G78gat), .B(G106gat), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n343_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n342_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n333_), .A2(new_n337_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n334_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT93), .A3(new_n338_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n364_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n367_), .A2(new_n368_), .A3(new_n366_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT100), .B(KEYINPUT0), .Z(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n332_), .A2(new_n294_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n323_), .A2(new_n288_), .A3(new_n331_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n288_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n393_), .B2(new_n389_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n384_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT33), .B(new_n384_), .C1(new_n392_), .C2(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G64gat), .B(G92gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT19), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT94), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n263_), .A2(KEYINPUT96), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n254_), .A2(new_n255_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n260_), .A2(new_n412_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT95), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n269_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n278_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n271_), .A2(new_n417_), .B1(new_n418_), .B2(new_n248_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n260_), .A2(new_n268_), .A3(KEYINPUT95), .A4(new_n261_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n422_), .A2(KEYINPUT97), .A3(new_n357_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT97), .B1(new_n422_), .B2(new_n357_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n280_), .B2(new_n357_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n409_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n422_), .A2(KEYINPUT98), .A3(new_n357_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n280_), .B2(new_n357_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT98), .B1(new_n422_), .B2(new_n357_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n408_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n406_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n424_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(KEYINPUT97), .A3(new_n357_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n427_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n409_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n434_), .A3(new_n405_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n393_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n388_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT101), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT101), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n388_), .A2(new_n447_), .A3(new_n385_), .A4(new_n391_), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n384_), .B(new_n444_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n400_), .A2(new_n443_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n392_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n384_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n394_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n396_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n431_), .B1(new_n357_), .B2(new_n422_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n408_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT32), .A3(new_n405_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n441_), .A2(KEYINPUT102), .A3(new_n434_), .A4(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n423_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n434_), .B(new_n459_), .C1(new_n461_), .C2(new_n409_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT102), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND4_X1   g263(.A1(new_n454_), .A2(new_n458_), .A3(new_n460_), .A4(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n306_), .B(new_n379_), .C1(new_n450_), .C2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n301_), .A2(new_n305_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n339_), .A2(new_n340_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n342_), .A2(new_n369_), .B1(new_n468_), .B2(new_n365_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n374_), .A2(new_n377_), .A3(new_n375_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n306_), .A2(new_n370_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n454_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT27), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n443_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT103), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n442_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n457_), .B2(new_n406_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n442_), .A2(new_n477_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .A4(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n247_), .B1(new_n466_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT104), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G190gat), .B(G218gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G134gat), .B(G162gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  NAND2_X1  g286(.A1(G232gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT34), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT35), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(KEYINPUT67), .A2(G85gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT67), .A2(G85gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(G92gat), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(G85gat), .B2(G92gat), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n499_), .A2(new_n500_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n501_), .A2(KEYINPUT68), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT65), .B(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n492_), .A2(KEYINPUT10), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT10), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G99gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT64), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT64), .B1(new_n508_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT66), .B(new_n507_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT71), .B1(G85gat), .B2(G92gat), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(G85gat), .B2(G92gat), .ZN(new_n519_));
  OAI221_X1 g318(.A(KEYINPUT69), .B1(KEYINPUT70), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT69), .B1(KEYINPUT70), .B2(KEYINPUT7), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n494_), .A2(new_n525_), .A3(new_n495_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(new_n519_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n517_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT72), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n517_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n490_), .B1(new_n536_), .B2(new_n223_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n489_), .A2(KEYINPUT35), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT76), .Z(new_n539_));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n540_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n517_), .A2(new_n531_), .A3(new_n222_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n537_), .A2(new_n542_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n517_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n534_), .B1(new_n517_), .B2(new_n531_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n223_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n490_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n543_), .A3(new_n544_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n541_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n487_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT77), .B1(new_n545_), .B2(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n487_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(KEYINPUT36), .A2(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n550_), .B(new_n542_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n556_), .B(new_n487_), .C1(new_n557_), .C2(KEYINPUT77), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT37), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(G231gat), .ZN(new_n564_));
  INV_X1    g363(.A(G233gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n219_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(G231gat), .B(G233gat), .C1(new_n216_), .C2(new_n218_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n569_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  INV_X1    g378(.A(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT16), .B(G183gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n566_), .A2(new_n575_), .A3(new_n567_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n577_), .A2(new_n578_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n578_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n577_), .A2(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n588_), .B2(KEYINPUT81), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT81), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n590_), .B(new_n586_), .C1(new_n577_), .C2(new_n584_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT82), .B(new_n585_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n584_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n575_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT81), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n586_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(KEYINPUT81), .A3(new_n587_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT82), .B1(new_n599_), .B2(new_n585_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n593_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n563_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n576_), .A2(KEYINPUT12), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n517_), .A2(new_n531_), .A3(new_n575_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n532_), .A2(new_n576_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n605_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n606_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT5), .B(G176gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT74), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT75), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n484_), .A2(new_n602_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(KEYINPUT105), .B2(KEYINPUT38), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G1gat), .A3(new_n474_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n601_), .A2(new_n559_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n636_), .A2(new_n627_), .A3(new_n483_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n207_), .B1(new_n637_), .B2(new_n454_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT106), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(G1324gat));
  NAND2_X1  g439(.A1(new_n481_), .A2(new_n476_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n208_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT39), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n208_), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n637_), .B2(new_n467_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n631_), .A2(new_n647_), .A3(new_n467_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n379_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n637_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n631_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n559_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n593_), .A2(new_n600_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n484_), .A2(new_n627_), .A3(new_n660_), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n661_), .A2(G29gat), .A3(new_n474_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n466_), .A2(new_n482_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n555_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n561_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT43), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n663_), .B(new_n668_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n670_), .A2(new_n627_), .A3(new_n601_), .A4(new_n246_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n454_), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT107), .B1(new_n675_), .B2(G29gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n662_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n641_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n661_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  INV_X1    g482(.A(new_n641_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n680_), .B1(new_n673_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT46), .ZN(G1329gat));
  XNOR2_X1  g487(.A(KEYINPUT108), .B(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n661_), .B2(new_n306_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n673_), .A2(G43gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n674_), .A2(new_n467_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g493(.A1(new_n661_), .A2(new_n379_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(G50gat), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n673_), .A2(G50gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n379_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(G1331gat));
  NOR4_X1   g498(.A1(new_n563_), .A2(new_n627_), .A3(new_n601_), .A4(new_n246_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n663_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n454_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n629_), .A2(new_n247_), .A3(new_n663_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n636_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n474_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(G57gat), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n708_), .A3(new_n641_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n705_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(new_n641_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n705_), .B2(new_n306_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n702_), .A2(new_n289_), .A3(new_n467_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  OR3_X1    g518(.A1(new_n701_), .A2(G78gat), .A3(new_n379_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G78gat), .B1(new_n705_), .B2(new_n379_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT50), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT50), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT110), .ZN(G1335gat));
  AND2_X1   g524(.A1(new_n704_), .A2(new_n660_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n454_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(G85gat), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n729_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n659_), .A2(new_n627_), .A3(new_n246_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n670_), .A2(new_n732_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n454_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n730_), .A2(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n726_), .B2(new_n641_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n641_), .A2(G92gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n733_), .B2(new_n737_), .ZN(G1337gat));
  AOI21_X1  g537(.A(new_n492_), .B1(new_n733_), .B2(new_n467_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n511_), .A2(new_n512_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n306_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n726_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1338gat));
  AOI21_X1  g543(.A(new_n668_), .B1(new_n563_), .B2(new_n663_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n669_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n653_), .B(new_n732_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT114), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n670_), .A2(new_n749_), .A3(new_n653_), .A4(new_n732_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(G106gat), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT115), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n748_), .A2(new_n753_), .A3(G106gat), .A4(new_n750_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(KEYINPUT52), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n726_), .A2(new_n507_), .A3(new_n653_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT113), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(KEYINPUT115), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n755_), .A2(new_n757_), .A3(new_n762_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(new_n471_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n641_), .A2(new_n474_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n604_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n613_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n604_), .A2(KEYINPUT55), .A3(new_n610_), .A4(new_n607_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n611_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n611_), .B2(new_n773_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n771_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n620_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n604_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n778_), .A2(KEYINPUT55), .B1(new_n768_), .B2(new_n613_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT117), .B1(new_n778_), .B2(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n611_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n621_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n777_), .A2(new_n623_), .A3(new_n246_), .A4(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n244_), .A2(new_n231_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n230_), .A2(new_n232_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n204_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n233_), .A2(new_n240_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n204_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n624_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n785_), .A2(new_n791_), .ZN(new_n792_));
  AND4_X1   g591(.A1(new_n767_), .A2(new_n792_), .A3(KEYINPUT57), .A4(new_n658_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n559_), .B1(new_n785_), .B2(new_n791_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n767_), .B1(new_n794_), .B2(KEYINPUT57), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n782_), .A2(new_n783_), .A3(new_n621_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n783_), .B1(new_n782_), .B2(new_n621_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n623_), .A4(new_n790_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n777_), .A2(new_n790_), .A3(new_n623_), .A4(new_n784_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n803_), .A3(new_n563_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n794_), .A2(KEYINPUT57), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n659_), .B1(new_n796_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n664_), .A2(new_n665_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n246_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n659_), .A4(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n560_), .A2(new_n659_), .A3(new_n810_), .A4(new_n562_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n813_), .A3(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n765_), .B(new_n766_), .C1(new_n807_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G113gat), .B1(new_n820_), .B2(new_n246_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n822_));
  INV_X1    g621(.A(new_n766_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n792_), .A2(KEYINPUT57), .A3(new_n658_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n792_), .A2(new_n658_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n800_), .A2(new_n803_), .A3(new_n563_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n794_), .A2(new_n767_), .A3(KEYINPUT57), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n825_), .A2(new_n828_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n601_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n811_), .A2(new_n813_), .A3(KEYINPUT54), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT54), .B1(new_n811_), .B2(new_n813_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n823_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n765_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n822_), .A2(new_n838_), .A3(new_n246_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n821_), .B1(new_n839_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n627_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n820_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n822_), .A2(new_n838_), .A3(new_n629_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n841_), .ZN(G1341gat));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  OAI21_X1  g645(.A(G127gat), .B1(new_n601_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT119), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n822_), .A2(new_n838_), .A3(new_n847_), .A4(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n819_), .B2(new_n601_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n808_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT120), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n822_), .A2(new_n838_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n819_), .B2(new_n658_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1343gat));
  INV_X1    g657(.A(new_n472_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n766_), .C1(new_n807_), .C2(new_n818_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n247_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n308_), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n630_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n309_), .ZN(G1345gat));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n860_), .B2(new_n601_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n836_), .A2(new_n867_), .A3(new_n659_), .A4(new_n859_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  INV_X1    g670(.A(G162gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n860_), .A2(new_n872_), .A3(new_n808_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n860_), .B2(new_n658_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT122), .B(new_n872_), .C1(new_n860_), .C2(new_n658_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n684_), .A2(new_n454_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n471_), .B(new_n880_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n246_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n765_), .B(new_n879_), .C1(new_n807_), .C2(new_n818_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884_), .B2(new_n247_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n883_), .B(new_n887_), .C1(new_n249_), .C2(new_n882_), .ZN(G1348gat));
  INV_X1    g687(.A(new_n627_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n881_), .B2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n881_), .A2(G176gat), .A3(new_n629_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT123), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n881_), .A2(new_n893_), .A3(G176gat), .A4(new_n629_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n892_), .B2(new_n894_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n884_), .A2(new_n601_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n271_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n258_), .B2(new_n896_), .ZN(G1350gat));
  AOI21_X1  g697(.A(new_n259_), .B1(new_n881_), .B2(new_n563_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n559_), .A2(new_n417_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n884_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT124), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G190gat), .B1(new_n884_), .B2(new_n808_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(new_n904_), .C1(new_n884_), .C2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1351gat));
  OAI211_X1 g705(.A(new_n859_), .B(new_n879_), .C1(new_n807_), .C2(new_n818_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n247_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n347_), .ZN(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n630_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n345_), .ZN(G1353gat));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n659_), .B1(new_n912_), .B2(new_n580_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n907_), .A2(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n914_), .B(new_n917_), .ZN(G1354gat));
  OAI21_X1  g717(.A(KEYINPUT127), .B1(new_n907_), .B2(new_n658_), .ZN(new_n919_));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n880_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(new_n559_), .A4(new_n859_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n919_), .A2(new_n920_), .A3(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n907_), .A2(new_n920_), .A3(new_n808_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1355gat));
endmodule


