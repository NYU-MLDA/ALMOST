//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(G169gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT26), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n222_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT83), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n210_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT91), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n231_), .A2(new_n232_), .A3(new_n237_), .A4(new_n234_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n230_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AOI211_X1 g040(.A(KEYINPUT92), .B(new_n230_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n219_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT21), .B(new_n244_), .C1(new_n245_), .C2(KEYINPUT87), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G197gat), .B(G204gat), .Z(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(KEYINPUT21), .B2(new_n245_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n246_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n243_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n231_), .A2(new_n232_), .A3(new_n215_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n218_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n233_), .B1(new_n213_), .B2(new_n211_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n227_), .B2(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n223_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n257_), .B(new_n222_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n263_), .B2(new_n253_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT90), .B(KEYINPUT20), .C1(new_n263_), .C2(new_n253_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n209_), .B1(new_n254_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n253_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n270_), .B(new_n219_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n253_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT20), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(new_n208_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n206_), .B1(new_n269_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n206_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n267_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n253_), .B2(new_n243_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n275_), .C1(new_n280_), .C2(new_n209_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(KEYINPUT94), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT94), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(new_n206_), .C1(new_n269_), .C2(new_n276_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n254_), .A2(new_n268_), .A3(new_n209_), .ZN(new_n287_));
  AOI211_X1 g086(.A(new_n253_), .B(new_n239_), .C1(new_n218_), .C2(new_n216_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n208_), .B1(new_n288_), .B2(new_n273_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n206_), .B(KEYINPUT97), .Z(new_n291_));
  OAI211_X1 g090(.A(KEYINPUT27), .B(new_n281_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  INV_X1    g093(.A(G141gat), .ZN(new_n295_));
  INV_X1    g094(.A(G148gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G141gat), .B(G148gat), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n304_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n253_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT89), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n253_), .B(new_n316_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n253_), .A2(KEYINPUT88), .ZN(new_n321_));
  INV_X1    g120(.A(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G228gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(KEYINPUT86), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(KEYINPUT86), .B2(new_n323_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n319_), .A3(new_n318_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G22gat), .B(G50gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n311_), .A2(KEYINPUT29), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n332_), .A2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n331_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n331_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n327_), .A2(new_n329_), .A3(new_n340_), .A4(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n293_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n311_), .A2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n305_), .B(new_n310_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n311_), .A2(new_n355_), .A3(new_n351_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT95), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n311_), .A2(KEYINPUT95), .A3(new_n355_), .A4(new_n351_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n364_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(new_n370_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT84), .B(G43gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n263_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(new_n351_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(G15gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT30), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT31), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n381_), .B(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n376_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n346_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT100), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n352_), .A2(new_n362_), .A3(new_n353_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n370_), .B(new_n391_), .C1(new_n360_), .C2(new_n362_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n373_), .A2(KEYINPUT33), .A3(new_n370_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n269_), .A2(new_n276_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n375_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n344_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT96), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n405_), .B(new_n344_), .C1(new_n397_), .C2(new_n402_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n376_), .A2(new_n344_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n286_), .A2(new_n407_), .A3(new_n292_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n286_), .A2(new_n407_), .A3(KEYINPUT98), .A4(new_n292_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n404_), .A2(new_n406_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n387_), .B(KEYINPUT85), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT99), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n390_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G229gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G1gat), .B(G8gat), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT77), .B(G15gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G22gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425_));
  INV_X1    g224(.A(G1gat), .ZN(new_n426_));
  INV_X1    g225(.A(G8gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT14), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n422_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(new_n428_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT78), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n421_), .A3(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G29gat), .B(G36gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT76), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n435_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n440_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AOI211_X1 g244(.A(KEYINPUT81), .B(new_n440_), .C1(new_n431_), .C2(new_n435_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n420_), .B(new_n441_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G113gat), .B(G141gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G169gat), .B(G197gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n440_), .A2(KEYINPUT15), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n440_), .A2(KEYINPUT15), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n443_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n445_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n446_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n447_), .B(new_n451_), .C1(new_n457_), .C2(new_n420_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n445_), .A2(new_n446_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n419_), .B1(new_n460_), .B2(new_n454_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n451_), .B1(new_n461_), .B2(new_n447_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G71gat), .B(G78gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(G57gat), .B(G64gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(KEYINPUT11), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT11), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n465_), .B2(KEYINPUT11), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT67), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n464_), .A4(new_n468_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n475_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT12), .B1(new_n479_), .B2(KEYINPUT71), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  AOI211_X1 g295(.A(KEYINPUT8), .B(new_n487_), .C1(new_n491_), .C2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n494_), .B1(G99gat), .B2(G106gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n488_), .B(new_n502_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n498_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT68), .B1(new_n497_), .B2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n493_), .A2(new_n495_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n488_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT8), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n498_), .A3(new_n506_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n501_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(KEYINPUT64), .A3(new_n501_), .A4(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n483_), .A2(KEYINPUT9), .ZN(new_n524_));
  AND2_X1   g323(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n484_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n527_), .A2(new_n496_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n523_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n523_), .B2(new_n529_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n516_), .A2(KEYINPUT70), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT70), .B1(new_n516_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n481_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n512_), .A2(new_n514_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n523_), .A2(new_n529_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n476_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n476_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n536_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n537_), .B1(new_n546_), .B2(new_n541_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT73), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(KEYINPUT74), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n556_), .A2(new_n558_), .A3(KEYINPUT13), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT13), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n452_), .A2(new_n453_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n540_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n569_));
  AOI22_X1  g368(.A1(new_n565_), .A2(new_n444_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(new_n572_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT36), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n578_), .B(KEYINPUT36), .Z(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT37), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n436_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n476_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n594_), .B1(new_n597_), .B2(new_n477_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n477_), .B2(new_n597_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n593_), .B(KEYINPUT17), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT80), .Z(new_n601_));
  OR2_X1    g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n588_), .A2(new_n604_), .ZN(new_n605_));
  NOR4_X1   g404(.A1(new_n418_), .A2(new_n463_), .A3(new_n562_), .A4(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n426_), .A3(new_n376_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n583_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n418_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n463_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n561_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n603_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n375_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n607_), .A2(new_n608_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  AOI21_X1  g418(.A(new_n427_), .B1(new_n615_), .B2(new_n293_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT39), .A3(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  INV_X1    g424(.A(new_n293_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(G8gat), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n624_), .A2(new_n625_), .B1(new_n606_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n628_), .A3(KEYINPUT40), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n616_), .B2(new_n413_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(KEYINPUT41), .A3(new_n636_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n413_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n606_), .A2(new_n383_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n344_), .B(KEYINPUT103), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n615_), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n606_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  NAND2_X1  g449(.A1(new_n603_), .A2(new_n610_), .ZN(new_n651_));
  NOR4_X1   g450(.A1(new_n418_), .A2(new_n463_), .A3(new_n562_), .A4(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n376_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n613_), .A2(new_n604_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n389_), .B(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n416_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n587_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n659_), .B2(new_n587_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n588_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n660_), .A3(new_n587_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n376_), .A2(G29gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n653_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT105), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n652_), .A2(new_n675_), .A3(new_n293_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n670_), .A2(new_n293_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n674_), .B(new_n678_), .C1(new_n679_), .C2(new_n675_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n670_), .B2(new_n293_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n678_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT105), .B(new_n673_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  INV_X1    g483(.A(G43gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n387_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n652_), .A2(new_n641_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT106), .B(G43gat), .Z(new_n688_));
  AOI22_X1  g487(.A1(new_n670_), .A2(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n652_), .A2(new_n692_), .A3(new_n646_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n665_), .A2(KEYINPUT107), .A3(new_n345_), .A4(new_n669_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n665_), .A2(new_n345_), .A3(new_n669_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n694_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  AND4_X1   g499(.A1(new_n694_), .A2(new_n699_), .A3(G50gat), .A4(new_n695_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n693_), .B1(new_n700_), .B2(new_n701_), .ZN(G1331gat));
  NOR3_X1   g501(.A1(new_n561_), .A2(new_n603_), .A3(new_n612_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n611_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n375_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n605_), .A2(new_n561_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n418_), .A3(new_n612_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n376_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n704_), .B2(new_n293_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n713_), .A3(new_n293_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n705_), .B2(new_n413_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n413_), .A2(G71gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT111), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n709_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n704_), .B2(new_n646_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT50), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n709_), .A2(new_n725_), .A3(new_n646_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1335gat));
  NOR4_X1   g528(.A1(new_n418_), .A2(new_n612_), .A3(new_n561_), .A4(new_n651_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G85gat), .B1(new_n730_), .B2(new_n376_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n562_), .A2(new_n463_), .A3(new_n603_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n376_), .B1(new_n526_), .B2(new_n525_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT112), .Z(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(new_n733_), .B2(new_n735_), .ZN(G1336gat));
  INV_X1    g535(.A(new_n733_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G92gat), .B1(new_n737_), .B2(new_n626_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n730_), .A2(new_n483_), .A3(new_n293_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n737_), .B2(new_n413_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n517_), .A2(new_n518_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n387_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n730_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n730_), .A2(new_n501_), .A3(new_n345_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n344_), .B(new_n732_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n501_), .B1(new_n749_), .B2(KEYINPUT113), .ZN(new_n750_));
  INV_X1    g549(.A(new_n732_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n345_), .B(new_n751_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n748_), .B1(new_n750_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G106gat), .B1(new_n752_), .B2(new_n753_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT113), .B1(new_n733_), .B2(new_n345_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(KEYINPUT52), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n747_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n747_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  INV_X1    g563(.A(new_n557_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n545_), .A2(KEYINPUT114), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n536_), .A2(new_n544_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(G230gat), .A3(G233gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n545_), .B2(KEYINPUT114), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT56), .B(new_n765_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n545_), .A2(KEYINPUT114), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n769_), .A3(new_n767_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n765_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n462_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n457_), .A2(new_n420_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n455_), .A2(new_n456_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n780_), .B(new_n451_), .C1(new_n420_), .C2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n549_), .A2(new_n555_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n779_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n764_), .B1(new_n778_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n785_), .A2(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT117), .A3(new_n772_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT58), .A3(new_n788_), .A4(new_n784_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n790_), .A2(new_n587_), .A3(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n556_), .A2(new_n558_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n779_), .A2(new_n782_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n785_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n556_), .B1(new_n458_), .B2(new_n779_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n785_), .B2(KEYINPUT115), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n583_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n583_), .A3(KEYINPUT116), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n794_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n603_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n588_), .A2(new_n463_), .A3(new_n561_), .A4(new_n604_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT54), .Z(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n387_), .A2(new_n375_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n346_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n612_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n810_), .B1(new_n807_), .B2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n795_), .A2(new_n796_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n783_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n776_), .B2(new_n765_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n829_), .B2(KEYINPUT56), .ZN(new_n830_));
  INV_X1    g629(.A(new_n801_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n804_), .B1(new_n832_), .B2(new_n610_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n808_), .A3(new_n806_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n790_), .A2(new_n587_), .A3(new_n793_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n824_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n603_), .B1(new_n825_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n815_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n839_), .A2(new_n840_), .B1(new_n820_), .B2(KEYINPUT59), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n841_), .A2(new_n612_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n823_), .B1(new_n842_), .B2(new_n822_), .ZN(G1340gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n562_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G120gat), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(G120gat), .B1(new_n562_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT119), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n846_), .B2(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n845_), .B1(new_n820_), .B2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n821_), .B2(new_n604_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n604_), .A2(G127gat), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT120), .Z(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n841_), .B2(new_n855_), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n841_), .A2(new_n587_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G134gat), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n583_), .A2(G134gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n820_), .B2(new_n859_), .ZN(G1343gat));
  AOI21_X1  g659(.A(new_n814_), .B1(new_n603_), .B2(new_n811_), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n641_), .A2(new_n375_), .A3(new_n293_), .A4(new_n344_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n612_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT121), .B(G141gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n562_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g668(.A1(new_n816_), .A2(new_n862_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT122), .B1(new_n870_), .B2(new_n603_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n864_), .A2(new_n872_), .A3(new_n604_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  NOR2_X1   g675(.A1(new_n870_), .A2(new_n583_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n587_), .A2(G162gat), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT123), .Z(new_n879_));
  OAI22_X1  g678(.A1(new_n877_), .A2(G162gat), .B1(new_n870_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1347gat));
  NOR3_X1   g681(.A1(new_n626_), .A2(new_n413_), .A3(new_n376_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n646_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n834_), .A2(new_n835_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n809_), .B1(new_n886_), .B2(KEYINPUT118), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n604_), .B1(new_n887_), .B2(new_n836_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n612_), .B(new_n885_), .C1(new_n888_), .C2(new_n814_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  OAI21_X1  g689(.A(G169gat), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n885_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n838_), .B2(new_n815_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT125), .B1(new_n893_), .B2(new_n612_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT62), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(KEYINPUT125), .A3(new_n612_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n889_), .A2(new_n890_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .A4(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n886_), .A2(KEYINPUT118), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n810_), .A3(new_n836_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n814_), .B1(new_n903_), .B2(new_n603_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n904_), .B2(new_n892_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT126), .B(new_n885_), .C1(new_n888_), .C2(new_n814_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT22), .B(G169gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n612_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n909_), .ZN(G1348gat));
  NOR2_X1   g709(.A1(new_n861_), .A2(new_n345_), .ZN(new_n911_));
  AND4_X1   g710(.A1(G176gat), .A2(new_n911_), .A3(new_n562_), .A4(new_n883_), .ZN(new_n912_));
  AOI21_X1  g711(.A(KEYINPUT126), .B1(new_n839_), .B2(new_n885_), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n901_), .B(new_n892_), .C1(new_n838_), .C2(new_n815_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n562_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(G176gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(KEYINPUT127), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n561_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(G176gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n912_), .B1(new_n917_), .B2(new_n920_), .ZN(G1349gat));
  NOR2_X1   g720(.A1(new_n884_), .A2(new_n603_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G183gat), .B1(new_n911_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n604_), .A2(new_n224_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n907_), .B2(new_n925_), .ZN(G1350gat));
  INV_X1    g725(.A(new_n907_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G190gat), .B1(new_n927_), .B2(new_n588_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n583_), .A2(new_n229_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1351gat));
  AND3_X1   g729(.A1(new_n413_), .A2(new_n293_), .A3(new_n407_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n816_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n612_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n562_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n604_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n932_), .B2(new_n588_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n583_), .A2(G218gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n932_), .B2(new_n944_), .ZN(G1355gat));
endmodule


