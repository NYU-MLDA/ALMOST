//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT68), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT68), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT68), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT8), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT9), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n221_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n212_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n221_), .A2(new_n230_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n206_), .A2(new_n209_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G232gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT34), .ZN(new_n236_));
  OAI22_X1  g035(.A1(new_n233_), .A2(new_n234_), .B1(KEYINPUT35), .B2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  OAI221_X1 g038(.A(new_n239_), .B1(KEYINPUT35), .B2(new_n236_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n236_), .A2(KEYINPUT35), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G190gat), .B(G218gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(G134gat), .B(G162gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(KEYINPUT36), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n240_), .B(new_n241_), .C1(new_n232_), .C2(new_n237_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT72), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT72), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n243_), .A2(new_n253_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n248_), .B(KEYINPUT36), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n243_), .B2(new_n250_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT37), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT37), .ZN(new_n260_));
  AOI211_X1 g059(.A(new_n260_), .B(new_n257_), .C1(new_n252_), .C2(new_n254_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G71gat), .B(G78gat), .Z(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(KEYINPUT11), .B2(new_n264_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n267_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n270_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT73), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n279_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G127gat), .B(G155gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT76), .ZN(new_n284_));
  XOR2_X1   g083(.A(G183gat), .B(G211gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT17), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n282_), .B(new_n290_), .C1(KEYINPUT17), .C2(new_n288_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n263_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n233_), .A2(new_n270_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT65), .B(KEYINPUT12), .Z(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n267_), .B(new_n269_), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n231_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G230gat), .A2(G233gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(KEYINPUT66), .A3(new_n303_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G120gat), .B(G148gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT5), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G176gat), .B(G204gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n310_), .A2(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT13), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n317_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n310_), .B(new_n315_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(new_n321_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n295_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT82), .B(G43gat), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332_));
  INV_X1    g131(.A(G169gat), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT81), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n333_), .A2(new_n334_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .A4(KEYINPUT24), .ZN(new_n346_));
  NOR2_X1   g145(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT80), .B(G183gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(KEYINPUT25), .ZN(new_n349_));
  INV_X1    g148(.A(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT26), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n340_), .B(new_n346_), .C1(new_n349_), .C2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(G190gat), .B2(new_n348_), .ZN(new_n359_));
  AND2_X1   g158(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n334_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n342_), .A2(new_n344_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(KEYINPUT30), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT30), .B1(new_n355_), .B2(new_n364_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n366_), .A2(G99gat), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G99gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n355_), .A2(new_n364_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n372_), .B2(new_n365_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n331_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G71gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(G99gat), .B1(new_n366_), .B2(new_n367_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n369_), .A3(new_n365_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n330_), .A3(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n374_), .B2(new_n381_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT31), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n381_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT31), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n382_), .A3(KEYINPUT83), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G127gat), .B(G134gat), .Z(new_n392_));
  XOR2_X1   g191(.A(G113gat), .B(G120gat), .Z(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G204gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G197gat), .ZN(new_n398_));
  INV_X1    g197(.A(G197gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(G204gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT21), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n397_), .B2(G197gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(G197gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n408_));
  OAI211_X1 g207(.A(new_n401_), .B(new_n402_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n407_), .A3(KEYINPUT21), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n370_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT19), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n338_), .B(new_n339_), .C1(G183gat), .C2(G190gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n363_), .A3(new_n362_), .ZN(new_n419_));
  AND2_X1   g218(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n351_), .B(new_n353_), .C1(new_n420_), .C2(new_n347_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n345_), .A2(KEYINPUT24), .A3(new_n341_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n421_), .A2(new_n358_), .A3(new_n422_), .A4(new_n335_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT20), .B1(new_n412_), .B2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n417_), .A2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G8gat), .B(G36gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT18), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n355_), .A2(new_n364_), .A3(new_n409_), .A4(new_n411_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n412_), .A2(new_n424_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT20), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n415_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n433_), .B2(new_n415_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n426_), .B(new_n430_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT27), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n412_), .C2(new_n424_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n413_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n415_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n433_), .A2(new_n415_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n430_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT99), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n442_), .B2(new_n415_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT99), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n430_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n438_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n426_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n447_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n437_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT27), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G141gat), .A2(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT2), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  NOR3_X1   g266(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n465_), .A2(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G141gat), .A2(G148gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n463_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n471_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n464_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n459_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT85), .B1(new_n459_), .B2(KEYINPUT1), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483_));
  INV_X1    g282(.A(G155gat), .ZN(new_n484_));
  INV_X1    g283(.A(G162gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT1), .ZN(new_n487_));
  AND2_X1   g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n486_), .A2(new_n460_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n479_), .B1(new_n482_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT87), .B1(new_n477_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n479_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n488_), .B2(new_n487_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n459_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n487_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n492_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n488_), .B1(new_n486_), .B2(new_n460_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n465_), .A2(new_n467_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n471_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n474_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n500_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n491_), .A2(KEYINPUT29), .A3(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n470_), .A2(new_n476_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n486_), .A2(new_n460_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n512_), .A2(new_n494_), .A3(new_n497_), .A4(new_n495_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n511_), .A2(new_n500_), .B1(new_n513_), .B2(new_n492_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n412_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n508_), .A2(new_n510_), .B1(new_n516_), .B2(new_n509_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n458_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n510_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n509_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT91), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G22gat), .B(G50gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n491_), .A2(new_n507_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n515_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n491_), .C2(new_n507_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n499_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n506_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n515_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT28), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n528_), .A2(new_n527_), .A3(new_n515_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n525_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n458_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n520_), .A2(new_n521_), .A3(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n522_), .A2(KEYINPUT91), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n517_), .A2(new_n518_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .A4(new_n458_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n524_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(KEYINPUT90), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n517_), .A2(new_n538_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n547_), .A2(new_n548_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n452_), .A2(new_n457_), .A3(new_n546_), .A4(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n394_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n491_), .A2(new_n507_), .A3(new_n394_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n395_), .A2(new_n514_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G225gat), .A2(G233gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT94), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n554_), .A2(new_n555_), .A3(new_n559_), .A4(new_n556_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n491_), .A2(new_n561_), .A3(new_n507_), .A4(new_n394_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n556_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT4), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n558_), .A2(new_n560_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G29gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G85gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT0), .B(G57gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n566_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR4_X1   g372(.A1(new_n396_), .A2(new_n552_), .A3(new_n553_), .A4(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n542_), .A2(new_n543_), .A3(new_n458_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n540_), .B1(new_n575_), .B2(KEYINPUT92), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n576_), .A2(new_n545_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(KEYINPUT33), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n558_), .A2(new_n560_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n554_), .A2(new_n555_), .A3(new_n563_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n454_), .A2(new_n581_), .A3(new_n437_), .A4(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n564_), .A2(new_n565_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n580_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n571_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n566_), .A2(new_n570_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n426_), .B(KEYINPUT96), .C1(new_n435_), .C2(new_n436_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n449_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n426_), .B(new_n597_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n594_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n591_), .A2(new_n592_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n577_), .B1(new_n588_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT98), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n546_), .A2(new_n551_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n603_), .A2(new_n457_), .A3(new_n452_), .A4(new_n572_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n577_), .B(new_n605_), .C1(new_n588_), .C2(new_n600_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n391_), .B(new_n395_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n574_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n212_), .A2(new_n278_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n210_), .A2(new_n278_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n234_), .A2(new_n277_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT78), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT78), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n613_), .B(new_n623_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(KEYINPUT79), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n609_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n329_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n272_), .A3(new_n573_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n630_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n326_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n255_), .A2(new_n258_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n637_), .A2(new_n609_), .A3(new_n294_), .A4(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n272_), .B1(new_n640_), .B2(new_n573_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n452_), .A2(new_n457_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n646_), .B2(G8gat), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT101), .B(new_n273_), .C1(new_n640_), .C2(new_n645_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(KEYINPUT39), .A3(new_n651_), .ZN(new_n652_));
  AND4_X1   g451(.A1(new_n273_), .A2(new_n329_), .A3(new_n645_), .A4(new_n631_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  NOR2_X1   g458(.A1(new_n396_), .A2(new_n553_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n376_), .B1(new_n640_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n632_), .A2(new_n376_), .A3(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n640_), .B2(new_n603_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n632_), .A2(new_n665_), .A3(new_n603_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n609_), .B2(new_n262_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n606_), .A2(new_n604_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n446_), .A2(new_n594_), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n674_), .A2(new_n593_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n572_), .A2(new_n675_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n605_), .B1(new_n676_), .B2(new_n577_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n608_), .B1(new_n673_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n552_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n660_), .A2(new_n679_), .A3(new_n572_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n263_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n672_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n326_), .A2(new_n636_), .A3(new_n294_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n688_), .B(new_n685_), .C1(new_n672_), .C2(new_n683_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n671_), .B1(new_n690_), .B2(new_n573_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n638_), .A2(new_n293_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n631_), .A2(new_n326_), .A3(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(new_n671_), .A3(new_n573_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n696_), .A3(new_n645_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT104), .B1(new_n690_), .B2(new_n645_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n682_), .B1(new_n681_), .B2(new_n263_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT43), .B(new_n262_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n686_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n688_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(KEYINPUT104), .A3(new_n645_), .A4(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT106), .B(new_n699_), .C1(new_n700_), .C2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n699_), .B1(new_n700_), .B2(new_n707_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT106), .B1(new_n711_), .B2(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT46), .B1(new_n708_), .B2(new_n709_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n714_), .A2(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT108), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n690_), .A2(G43gat), .A3(new_n660_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n693_), .A2(new_n660_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(G43gat), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n693_), .B2(new_n603_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n603_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n690_), .B2(new_n727_), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n609_), .A2(new_n639_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n326_), .A2(new_n636_), .A3(new_n294_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n572_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n609_), .A2(new_n636_), .A3(new_n326_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n295_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n573_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n731_), .B2(new_n645_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT48), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n739_), .A3(new_n645_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n731_), .B2(new_n660_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT49), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n735_), .A2(new_n744_), .A3(new_n660_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT109), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n731_), .B2(new_n603_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n735_), .A2(new_n750_), .A3(new_n603_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  AND2_X1   g554(.A1(new_n734_), .A2(new_n692_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n222_), .A3(new_n573_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n326_), .A2(new_n636_), .A3(new_n293_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n684_), .A2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n573_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(new_n222_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n223_), .A3(new_n645_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n645_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n223_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n660_), .A3(new_n226_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT111), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n369_), .B1(new_n759_), .B2(new_n660_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g569(.A(new_n227_), .B1(new_n759_), .B2(new_n603_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n227_), .A3(new_n603_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g576(.A1(new_n306_), .A2(new_n307_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n300_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n308_), .A2(KEYINPUT55), .ZN(new_n783_));
  INV_X1    g582(.A(new_n302_), .ZN(new_n784_));
  OAI211_X1 g583(.A(G230gat), .B(G233gat), .C1(new_n300_), .C2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n314_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n314_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(KEYINPUT114), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n314_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT114), .A3(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n628_), .A2(new_n316_), .A3(new_n629_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n789_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n788_), .B2(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n791_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n314_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n797_), .B(new_n798_), .C1(new_n801_), .C2(KEYINPUT114), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n623_), .B1(new_n615_), .B2(new_n612_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n323_), .A2(new_n627_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n796_), .A2(new_n802_), .A3(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n638_), .A3(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n316_), .A2(new_n627_), .A3(new_n805_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n262_), .B1(new_n812_), .B2(KEYINPUT58), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(KEYINPUT58), .B2(new_n812_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n809_), .B1(new_n807_), .B2(new_n638_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n294_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n327_), .B2(new_n636_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n295_), .A2(new_n819_), .A3(new_n630_), .A4(new_n326_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n660_), .A2(new_n679_), .A3(new_n573_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT117), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G113gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n636_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT59), .B1(new_n822_), .B2(KEYINPUT118), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n825_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n822_), .B(new_n824_), .C1(KEYINPUT118), .C2(KEYINPUT59), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n630_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n827_), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n326_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n826_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n326_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n839_), .A3(new_n293_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n294_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n826_), .A2(new_n843_), .A3(new_n639_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n262_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n843_), .ZN(G1343gat));
  NOR4_X1   g645(.A1(new_n660_), .A2(new_n577_), .A3(new_n645_), .A4(new_n572_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT119), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n822_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n630_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT120), .B(G141gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n326_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT121), .B(G148gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1345gat));
  NOR2_X1   g654(.A1(new_n849_), .A2(new_n294_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  OAI21_X1  g657(.A(G162gat), .B1(new_n849_), .B2(new_n262_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n639_), .A2(new_n485_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n849_), .B2(new_n860_), .ZN(G1347gat));
  NAND3_X1  g660(.A1(new_n660_), .A2(new_n645_), .A3(new_n572_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT122), .Z(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n603_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n822_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI211_X1 g665(.A(KEYINPUT62), .B(new_n333_), .C1(new_n866_), .C2(new_n636_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n636_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G169gat), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n866_), .B(new_n636_), .C1(new_n361_), .C2(new_n360_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(G1348gat));
  NOR2_X1   g671(.A1(new_n865_), .A2(new_n326_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n334_), .ZN(G1349gat));
  OAI21_X1  g673(.A(new_n348_), .B1(new_n865_), .B2(new_n294_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n420_), .A2(new_n347_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n865_), .A2(new_n877_), .A3(new_n294_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT123), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n866_), .A2(new_n293_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n880_), .B(new_n875_), .C1(new_n881_), .C2(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n865_), .B2(new_n262_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n638_), .A2(new_n354_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n865_), .B2(new_n885_), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n807_), .A2(new_n638_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n808_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n814_), .A3(new_n810_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n889_), .A2(new_n294_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n608_), .A2(new_n603_), .A3(new_n645_), .A4(new_n572_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT124), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  INV_X1    g692(.A(new_n891_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n822_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n630_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n399_), .ZN(G1352gat));
  AOI21_X1  g696(.A(new_n326_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT125), .B(G204gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n893_), .B1(new_n822_), .B2(new_n894_), .ZN(new_n901_));
  AOI211_X1 g700(.A(KEYINPUT124), .B(new_n891_), .C1(new_n817_), .C2(new_n821_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n293_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT63), .B(G211gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n294_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n903_), .A2(KEYINPUT126), .A3(new_n908_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n905_), .B1(new_n910_), .B2(new_n911_), .ZN(G1354gat));
  NAND2_X1  g711(.A1(new_n892_), .A2(new_n895_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n639_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT127), .B(G218gat), .Z(new_n915_));
  NOR2_X1   g714(.A1(new_n262_), .A2(new_n915_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n915_), .B1(new_n913_), .B2(new_n916_), .ZN(G1355gat));
endmodule


