//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(G15gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT22), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT79), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT80), .B(G176gat), .Z(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(KEYINPUT22), .B2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT23), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT74), .B(G190gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(G183gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229_));
  OAI21_X1  g028(.A(G190gat), .B1(new_n229_), .B2(KEYINPUT26), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT75), .ZN(new_n232_));
  OAI221_X1 g031(.A(new_n228_), .B1(new_n230_), .B2(new_n232_), .C1(new_n220_), .C2(new_n231_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n218_), .A2(new_n215_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n215_), .A2(KEYINPUT23), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n227_), .B(new_n233_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  OAI22_X1  g039(.A1(new_n214_), .A2(new_n224_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n241_), .A2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n206_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n241_), .A2(new_n244_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n205_), .A3(new_n245_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT31), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G127gat), .B(G134gat), .Z(new_n257_));
  XOR2_X1   g056(.A(G113gat), .B(G120gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n248_), .A2(new_n250_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n251_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT31), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n253_), .A3(new_n264_), .A4(new_n252_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n256_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n260_), .B1(new_n256_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  XOR2_X1   g070(.A(G197gat), .B(G204gat), .Z(new_n272_));
  XOR2_X1   g071(.A(G211gat), .B(G218gat), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(KEYINPUT21), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G204gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(KEYINPUT21), .B(new_n280_), .C1(new_n272_), .C2(KEYINPUT84), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n281_), .A3(KEYINPUT85), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n275_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n235_), .A2(new_n236_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n223_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT22), .B(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n292_), .B2(new_n211_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n226_), .A2(new_n223_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n228_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n225_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n300_), .A2(new_n219_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT90), .Z(new_n305_));
  AOI21_X1  g104(.A(new_n286_), .B1(new_n297_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n284_), .A2(new_n285_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n274_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT20), .B1(new_n308_), .B2(new_n241_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n271_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n297_), .A2(new_n305_), .A3(new_n286_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n271_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n308_), .B2(new_n241_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G64gat), .B(G92gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n310_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(KEYINPUT27), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n308_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n286_), .A2(KEYINPUT86), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n327_), .A2(new_n297_), .A3(new_n328_), .A4(new_n304_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n312_), .B1(new_n329_), .B2(new_n314_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n306_), .A2(new_n309_), .A3(new_n271_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n321_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n269_), .A2(new_n324_), .B1(new_n325_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n339_), .B(KEYINPUT3), .Z(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT2), .Z(new_n342_));
  OAI211_X1 g141(.A(new_n336_), .B(new_n338_), .C1(new_n340_), .C2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n337_), .B1(KEYINPUT1), .B2(new_n336_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(KEYINPUT1), .B2(new_n336_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n260_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n335_), .B1(new_n349_), .B2(KEYINPUT4), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT93), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n343_), .A2(new_n259_), .A3(new_n347_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT93), .B1(new_n356_), .B2(new_n350_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n353_), .A3(new_n334_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT95), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n349_), .A2(new_n360_), .A3(new_n353_), .A4(new_n334_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n357_), .A3(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n355_), .A2(new_n357_), .A3(new_n362_), .A4(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n348_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT83), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n308_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n375_), .B(new_n382_), .C1(new_n383_), .C2(new_n380_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n286_), .A2(KEYINPUT86), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n326_), .B(new_n275_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n380_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n375_), .B1(new_n390_), .B2(new_n382_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT88), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n382_), .B1(new_n383_), .B2(new_n380_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n374_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n384_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n377_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G22gat), .B(G50gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n384_), .B2(KEYINPUT87), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n333_), .B(new_n373_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n372_), .B(new_n408_), .C1(new_n316_), .C2(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n371_), .A2(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n354_), .B(new_n334_), .C1(KEYINPUT4), .C2(new_n349_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n349_), .A2(new_n353_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n368_), .B1(new_n413_), .B2(new_n335_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n371_), .A2(new_n410_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(new_n415_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n385_), .A2(new_n391_), .A3(KEYINPUT88), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n395_), .B1(new_n394_), .B2(new_n384_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n384_), .A2(KEYINPUT87), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n418_), .A2(new_n419_), .B1(new_n420_), .B2(new_n401_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n403_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n268_), .B1(new_n406_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n256_), .A2(new_n265_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n259_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n256_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n373_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n333_), .A2(new_n403_), .A3(new_n421_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(G85gat), .A2(G92gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  INV_X1    g239(.A(G106gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n433_), .B1(new_n438_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n435_), .A2(new_n437_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n443_), .A3(new_n442_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n446_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n433_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT9), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n448_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT10), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n440_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n441_), .A3(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n455_), .A2(KEYINPUT9), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n457_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n433_), .A2(KEYINPUT9), .B1(new_n435_), .B2(new_n437_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n455_), .A2(KEYINPUT9), .ZN(new_n467_));
  AND2_X1   g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n470_), .B2(new_n441_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT64), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n447_), .B(new_n451_), .C1(new_n465_), .C2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G29gat), .B(G36gat), .Z(new_n474_));
  XOR2_X1   g273(.A(G43gat), .B(G50gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G232gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT34), .ZN(new_n484_));
  INV_X1    g283(.A(new_n480_), .ZN(new_n485_));
  OAI221_X1 g284(.A(new_n482_), .B1(KEYINPUT35), .B2(new_n484_), .C1(new_n473_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(KEYINPUT35), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT69), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G190gat), .B(G218gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G134gat), .B(G162gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT36), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n489_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(KEYINPUT36), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n488_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499_));
  INV_X1    g298(.A(G8gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G71gat), .B(G78gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(KEYINPUT11), .ZN(new_n509_));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510_));
  INV_X1    g309(.A(G64gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G57gat), .ZN(new_n512_));
  INV_X1    g311(.A(G57gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G64gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n514_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n509_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n520_), .B(new_n509_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n506_), .B(new_n522_), .Z(new_n523_));
  XOR2_X1   g322(.A(G127gat), .B(G155gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT16), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G183gat), .B(G211gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  OR3_X1    g329(.A1(new_n523_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n506_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(new_n518_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n518_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n430_), .A2(new_n498_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n473_), .A2(new_n522_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n454_), .A2(new_n455_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n443_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n542_), .B(new_n446_), .C1(new_n545_), .C2(new_n448_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n450_), .B1(new_n449_), .B2(new_n433_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n464_), .B1(new_n457_), .B2(new_n463_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n466_), .A2(new_n471_), .A3(KEYINPUT64), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n548_), .A2(new_n521_), .A3(new_n519_), .A4(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n540_), .B1(new_n541_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT12), .B(new_n509_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n549_), .A2(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n447_), .A2(new_n451_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n548_), .A2(new_n551_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n552_), .B(new_n559_), .C1(new_n560_), .C2(KEYINPUT12), .ZN(new_n561_));
  INV_X1    g360(.A(new_n540_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n554_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n559_), .A2(new_n552_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT12), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n541_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n564_), .A2(KEYINPUT67), .A3(new_n540_), .A4(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n553_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G120gat), .B(G148gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n573_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n575_), .B(new_n576_), .C1(KEYINPUT68), .C2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n579_));
  INV_X1    g378(.A(new_n576_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n481_), .A2(new_n504_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n504_), .A2(new_n485_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n504_), .B(new_n485_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(G229gat), .A3(G233gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G113gat), .B(G141gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(KEYINPUT73), .A3(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n594_), .B1(new_n590_), .B2(KEYINPUT72), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(KEYINPUT72), .B2(new_n590_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n583_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n539_), .A2(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT97), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT97), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n202_), .B1(new_n608_), .B2(new_n372_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT98), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n430_), .A2(new_n603_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n498_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n495_), .A2(new_n497_), .A3(new_n612_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n538_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n582_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  AOI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(KEYINPUT96), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n372_), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(KEYINPUT96), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n610_), .A2(new_n623_), .ZN(G1324gat));
  INV_X1    g423(.A(new_n333_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n500_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n605_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n500_), .B1(new_n627_), .B2(new_n625_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n628_), .A2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n626_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n633_), .B(new_n635_), .ZN(G1325gat));
  NAND2_X1  g435(.A1(new_n608_), .A2(new_n268_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(G15gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n268_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n641_), .B2(new_n204_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n639_), .A2(KEYINPUT41), .A3(new_n642_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n618_), .A2(new_n204_), .A3(new_n268_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n421_), .A2(new_n403_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n608_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n618_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n498_), .A2(new_n538_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT104), .Z(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n583_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n611_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n659_), .A2(G29gat), .A3(new_n373_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n538_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n583_), .A2(new_n661_), .A3(new_n603_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n615_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n612_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n423_), .B2(new_n429_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT43), .B1(new_n666_), .B2(KEYINPUT101), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n662_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n662_), .B(KEYINPUT44), .C1(new_n667_), .C2(new_n668_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n372_), .A4(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(G29gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n372_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  AND4_X1   g477(.A1(KEYINPUT103), .A2(new_n677_), .A3(G29gat), .A4(new_n674_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n660_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n671_), .A2(new_n625_), .A3(new_n673_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n333_), .A2(G36gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n659_), .A2(KEYINPUT45), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT45), .B1(new_n659_), .B2(new_n685_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1329gat));
  AND2_X1   g490(.A1(new_n671_), .A2(new_n673_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(G43gat), .A3(new_n268_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n243_), .B1(new_n659_), .B2(new_n640_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(KEYINPUT47), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT47), .B1(new_n693_), .B2(new_n694_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1330gat));
  INV_X1    g496(.A(new_n650_), .ZN(new_n698_));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n658_), .A2(new_n650_), .A3(new_n611_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n692_), .A2(new_n700_), .B1(new_n699_), .B2(new_n701_), .ZN(G1331gat));
  NAND3_X1  g501(.A1(new_n539_), .A2(new_n583_), .A3(new_n603_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n373_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n430_), .A2(new_n602_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT106), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n665_), .A2(new_n582_), .A3(new_n538_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n372_), .A2(new_n513_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n704_), .B1(new_n708_), .B2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n703_), .B2(new_n333_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n625_), .A2(new_n511_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n708_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n703_), .B2(new_n640_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n640_), .A2(G71gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n708_), .B2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n703_), .B2(new_n698_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n698_), .A2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n708_), .B2(new_n721_), .ZN(G1335gat));
  OR2_X1    g521(.A1(new_n667_), .A2(new_n668_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n661_), .A2(new_n582_), .A3(new_n602_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n372_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G85gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n657_), .A2(new_n582_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n706_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n372_), .A2(new_n452_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1336gat));
  OAI21_X1  g530(.A(new_n453_), .B1(new_n729_), .B2(new_n333_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n333_), .A2(new_n453_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n734_), .A2(new_n735_), .B1(new_n725_), .B2(new_n736_), .ZN(G1337gat));
  INV_X1    g536(.A(new_n470_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n729_), .A2(new_n738_), .A3(new_n640_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n725_), .A2(new_n268_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G99gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(G1338gat));
  OAI211_X1 g542(.A(new_n650_), .B(new_n724_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G106gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G106gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n650_), .A2(new_n441_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n746_), .A2(new_n747_), .B1(new_n729_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g549(.A1(new_n640_), .A2(new_n373_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n428_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n584_), .A2(new_n586_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n585_), .B1(new_n754_), .B2(KEYINPUT113), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(KEYINPUT113), .B2(new_n754_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n594_), .B1(new_n588_), .B2(new_n585_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n599_), .A2(new_n576_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n559_), .A2(new_n552_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT12), .B1(new_n473_), .B2(new_n522_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT67), .B1(new_n765_), .B2(new_n540_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n561_), .A2(new_n554_), .A3(new_n562_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n762_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n562_), .A2(KEYINPUT55), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n566_), .A2(new_n552_), .A3(new_n559_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n562_), .A2(KEYINPUT110), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n561_), .B2(new_n771_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n760_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n761_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n763_), .A2(new_n764_), .A3(new_n771_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n771_), .B2(new_n770_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n775_), .A2(new_n777_), .A3(KEYINPUT111), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n572_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n768_), .A2(new_n773_), .A3(new_n760_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT111), .B1(new_n775_), .B2(new_n777_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n572_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n759_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT58), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n759_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n572_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n780_), .B(new_n573_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT114), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n788_), .A2(new_n665_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n788_), .A2(new_n665_), .A3(KEYINPUT115), .A4(new_n794_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n599_), .A2(new_n758_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n781_), .A2(KEYINPUT112), .A3(new_n785_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n602_), .A2(new_n576_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n791_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n801_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n799_), .B1(new_n806_), .B2(new_n498_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n498_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n802_), .A2(new_n805_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n808_), .C1(new_n809_), .C2(new_n801_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n797_), .A2(new_n798_), .A3(new_n807_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n538_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n616_), .A2(new_n582_), .A3(new_n603_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n753_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n602_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n816_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n810_), .A2(new_n795_), .A3(new_n807_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(new_n820_), .B2(new_n661_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  INV_X1    g621(.A(new_n753_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n602_), .B2(KEYINPUT116), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(KEYINPUT116), .B2(new_n826_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n817_), .B1(new_n825_), .B2(new_n828_), .ZN(G1340gat));
  OAI211_X1 g628(.A(new_n583_), .B(new_n824_), .C1(new_n816_), .C2(new_n822_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G120gat), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n816_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n832_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n837_), .A3(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n818_), .B2(new_n538_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n841_), .A2(KEYINPUT118), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(KEYINPUT118), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n661_), .A2(G127gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n842_), .A2(new_n843_), .B1(new_n825_), .B2(new_n845_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n816_), .B2(new_n498_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n665_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT119), .B(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT120), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n825_), .B2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n812_), .A2(new_n815_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n698_), .A2(new_n268_), .A3(new_n625_), .A4(new_n373_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n602_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g657(.A1(new_n855_), .A2(new_n582_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(G148gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n855_), .A2(new_n538_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OR3_X1    g663(.A1(new_n855_), .A2(G162gat), .A3(new_n808_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G162gat), .B1(new_n855_), .B2(new_n848_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1347gat));
  NAND3_X1  g666(.A1(new_n268_), .A2(new_n373_), .A3(new_n625_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n650_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n821_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870_), .B2(new_n603_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n873_));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n602_), .A3(new_n292_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n873_), .B2(new_n875_), .ZN(G1348gat));
  INV_X1    g675(.A(new_n211_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(new_n583_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n853_), .A2(new_n698_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(G176gat), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n868_), .A2(new_n582_), .A3(new_n884_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n880_), .A2(new_n881_), .B1(new_n883_), .B2(new_n885_), .ZN(G1349gat));
  NOR3_X1   g685(.A1(new_n870_), .A2(new_n228_), .A3(new_n538_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n868_), .A2(new_n538_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(G183gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n870_), .B2(new_n848_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT124), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n874_), .A2(new_n301_), .A3(new_n498_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  NOR4_X1   g694(.A1(new_n698_), .A2(new_n268_), .A3(new_n372_), .A4(new_n333_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n853_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n602_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n853_), .A2(new_n896_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n582_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n279_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n897_), .B2(new_n661_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  NOR3_X1   g704(.A1(new_n900_), .A2(new_n538_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n905_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n897_), .A2(new_n661_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n900_), .A2(new_n538_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n909_), .B(new_n910_), .C1(new_n911_), .C2(new_n903_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n907_), .A2(new_n912_), .ZN(G1354gat));
  XNOR2_X1  g712(.A(KEYINPUT126), .B(G218gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n900_), .A2(new_n848_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n897_), .A2(new_n498_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(G1355gat));
endmodule


