//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT80), .B(G15gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT77), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT76), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT76), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT25), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n210_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n207_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT76), .B(G183gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n216_), .B1(new_n226_), .B2(KEYINPUT25), .ZN(new_n227_));
  OAI211_X1 g026(.A(KEYINPUT77), .B(new_n223_), .C1(new_n227_), .C2(new_n210_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT23), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n221_), .A2(KEYINPUT24), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n225_), .A2(new_n228_), .A3(new_n233_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n230_), .A2(KEYINPUT79), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n232_), .A3(KEYINPUT79), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n238_), .B(new_n239_), .C1(G190gat), .C2(new_n226_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT78), .B(G169gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n236_), .A2(new_n237_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n237_), .B1(new_n236_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(G43gat), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT30), .ZN(new_n249_));
  INV_X1    g048(.A(G43gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n236_), .A2(new_n237_), .A3(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G99gat), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n247_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n206_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n245_), .A2(new_n246_), .A3(G43gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n250_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n247_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n205_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT31), .ZN(new_n265_));
  INV_X1    g064(.A(G120gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(G127gat), .A2(G134gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G127gat), .A2(G134gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT81), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT81), .B1(new_n267_), .B2(new_n268_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n270_), .A2(G113gat), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G113gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n276_), .B2(new_n269_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n266_), .B1(new_n272_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(G113gat), .B1(new_n270_), .B2(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n273_), .A3(new_n269_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(G120gat), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .A4(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n265_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n265_), .B2(new_n285_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n202_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n265_), .A2(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n265_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT83), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n296_));
  INV_X1    g095(.A(G155gat), .ZN(new_n297_));
  INV_X1    g096(.A(G162gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n301_), .B(new_n302_), .C1(new_n305_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(KEYINPUT1), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G155gat), .A3(G162gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n299_), .A2(new_n310_), .A3(new_n312_), .A4(new_n300_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(KEYINPUT85), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT85), .B1(new_n313_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n309_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n309_), .B(KEYINPUT86), .C1(new_n315_), .C2(new_n316_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n295_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G228gat), .ZN(new_n322_));
  INV_X1    g121(.A(G233gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G204gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G197gat), .ZN(new_n326_));
  INV_X1    g125(.A(G197gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G204gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT87), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n329_), .A2(KEYINPUT21), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT21), .B1(new_n329_), .B2(new_n330_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n328_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(new_n330_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n331_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n321_), .A2(new_n324_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n324_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n317_), .A2(KEYINPUT29), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n340_));
  OAI21_X1  g139(.A(G78gat), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n316_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n313_), .A2(KEYINPUT85), .A3(new_n314_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT86), .B1(new_n344_), .B2(new_n309_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n320_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT29), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n338_), .A3(new_n335_), .ZN(new_n348_));
  INV_X1    g147(.A(G78gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n340_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n341_), .A2(G106gat), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(G106gat), .B1(new_n341_), .B2(new_n351_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n294_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n319_), .A2(new_n295_), .A3(new_n320_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT28), .B(G22gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G50gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n355_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G106gat), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n337_), .A2(G78gat), .A3(new_n340_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n349_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n341_), .A2(G106gat), .A3(new_n351_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT88), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n294_), .B(new_n358_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n282_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n282_), .A2(new_n317_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n319_), .A2(new_n320_), .B1(new_n281_), .B2(new_n278_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(KEYINPUT4), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n282_), .A2(new_n317_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n374_), .A2(new_n377_), .A3(new_n369_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT91), .B(KEYINPUT0), .Z(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n387_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n376_), .A2(new_n379_), .A3(new_n384_), .A4(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n368_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n384_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n371_), .A2(new_n372_), .A3(new_n369_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT19), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n336_), .B1(new_n236_), .B2(new_n244_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n220_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n222_), .A3(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n216_), .A2(new_n403_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n238_), .A2(new_n404_), .A3(new_n239_), .A4(new_n223_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n405_), .B2(new_n234_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n406_), .B2(new_n335_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n397_), .B1(new_n398_), .B2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n409_));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n236_), .A2(new_n336_), .A3(new_n244_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n406_), .B2(new_n335_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n396_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n408_), .A2(new_n417_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n413_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n408_), .A2(KEYINPUT90), .A3(new_n413_), .A4(new_n417_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n388_), .A2(new_n390_), .A3(new_n394_), .A4(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT4), .B1(new_n374_), .B2(new_n377_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n371_), .A2(new_n370_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n368_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n392_), .B1(new_n430_), .B2(new_n378_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n385_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT93), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n421_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n396_), .B1(new_n398_), .B2(new_n407_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n414_), .A2(new_n397_), .A3(new_n416_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT94), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(KEYINPUT94), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n432_), .A2(new_n435_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n366_), .A2(new_n367_), .B1(new_n427_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n385_), .A2(new_n431_), .A3(KEYINPUT95), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT95), .B1(new_n385_), .B2(new_n431_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n446_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n425_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT97), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n438_), .A2(new_n413_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n423_), .A3(KEYINPUT27), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT96), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n423_), .A3(KEYINPUT96), .A4(KEYINPUT27), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n425_), .A2(KEYINPUT97), .A3(new_n448_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n443_), .B1(new_n447_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n293_), .A2(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n425_), .A2(KEYINPUT97), .A3(new_n448_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT97), .B1(new_n425_), .B2(new_n448_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT98), .B1(new_n465_), .B2(new_n457_), .ZN(new_n466_));
  AND4_X1   g265(.A1(KEYINPUT98), .A2(new_n451_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n290_), .A2(new_n291_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n366_), .A2(new_n367_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n468_), .A2(new_n446_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(KEYINPUT99), .A3(new_n468_), .A4(new_n446_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n462_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT10), .B(G99gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT64), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT65), .B(G106gat), .Z(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT66), .B(G92gat), .Z(new_n482_));
  INV_X1    g281(.A(G85gat), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n482_), .A2(KEYINPUT9), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G85gat), .B(G92gat), .Z(new_n485_));
  AND2_X1   g284(.A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT6), .Z(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n481_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  OR3_X1    g289(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT8), .B1(new_n485_), .B2(KEYINPUT67), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n490_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT11), .ZN(new_n505_));
  XOR2_X1   g304(.A(G57gat), .B(G64gat), .Z(new_n506_));
  OR3_X1    g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n505_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(KEYINPUT12), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n498_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n490_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n510_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n490_), .A2(new_n512_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n510_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .A4(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n514_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G176gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n325_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(new_n524_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(KEYINPUT69), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n534_), .A3(new_n529_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n535_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G29gat), .B(G36gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n250_), .ZN(new_n541_));
  INV_X1    g340(.A(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT15), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT74), .B(G8gat), .ZN(new_n545_));
  INV_X1    g344(.A(G1gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G8gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(G1gat), .ZN(new_n552_));
  INV_X1    g351(.A(G8gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n544_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT75), .Z(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n556_), .A2(new_n543_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n562_), .B2(new_n557_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n219_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n327_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n561_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n539_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n477_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G134gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n298_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n502_), .A2(new_n544_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n518_), .A2(new_n543_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT70), .Z(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT34), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT35), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n502_), .A2(new_n544_), .B1(new_n518_), .B2(new_n543_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(KEYINPUT71), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT71), .B1(new_n586_), .B2(new_n584_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n574_), .B(new_n578_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n589_), .B2(KEYINPUT71), .ZN(new_n593_));
  INV_X1    g392(.A(new_n577_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n578_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT73), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(KEYINPUT72), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n578_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n604_), .A3(new_n595_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT37), .A4(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n510_), .B(new_n608_), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n556_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n211_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(G211gat), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n610_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n616_), .B2(new_n610_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n607_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n573_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n446_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n546_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT38), .ZN(new_n625_));
  INV_X1    g424(.A(new_n599_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n573_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n446_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(G1324gat));
  OAI21_X1  g429(.A(G8gat), .B1(new_n628_), .B2(new_n468_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT39), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n465_), .A2(KEYINPUT98), .A3(new_n457_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n459_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n622_), .A2(new_n545_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT100), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n632_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1325gat));
  INV_X1    g441(.A(new_n293_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G15gat), .B1(new_n628_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n647_), .A3(new_n293_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1326gat));
  OAI21_X1  g448(.A(G22gat), .B1(new_n628_), .B2(new_n470_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT42), .ZN(new_n651_));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n470_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n622_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(new_n607_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n657_), .B(new_n658_), .C1(new_n477_), .C2(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n293_), .A2(new_n461_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n474_), .A2(new_n636_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT99), .B1(new_n662_), .B2(new_n446_), .ZN(new_n663_));
  NOR4_X1   g462(.A1(new_n474_), .A2(new_n636_), .A3(new_n472_), .A4(new_n623_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n657_), .A2(new_n658_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n665_), .A2(new_n607_), .A3(new_n666_), .A4(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n660_), .A2(new_n668_), .A3(new_n571_), .A4(new_n620_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n656_), .B1(new_n674_), .B2(new_n446_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT104), .B(new_n623_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(G29gat), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n599_), .A2(new_n619_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n573_), .A2(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n446_), .A2(G29gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n636_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G36gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n679_), .ZN(new_n685_));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n685_), .A2(KEYINPUT45), .A3(new_n686_), .A4(new_n636_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n573_), .A2(new_n686_), .A3(new_n678_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n468_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n682_), .B1(new_n684_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n682_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n694_), .B(new_n691_), .C1(new_n683_), .C2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1329gat));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n469_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G43gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n679_), .A2(G43gat), .A3(new_n643_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT47), .B(new_n700_), .C1(new_n698_), .C2(G43gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1330gat));
  OAI21_X1  g503(.A(G50gat), .B1(new_n674_), .B2(new_n470_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n685_), .A2(new_n542_), .A3(new_n653_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n477_), .A2(new_n569_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n539_), .A3(new_n627_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n446_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n708_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n539_), .A3(new_n621_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n714_), .A2(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(KEYINPUT107), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n623_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n711_), .B1(new_n717_), .B2(new_n710_), .ZN(G1332gat));
  NOR3_X1   g517(.A1(new_n714_), .A2(G64gat), .A3(new_n468_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G64gat), .B1(new_n709_), .B2(new_n468_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n709_), .B2(new_n643_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(G71gat), .C1(new_n709_), .C2(new_n643_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n643_), .A2(G71gat), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n725_), .A2(new_n728_), .B1(new_n714_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n709_), .B2(new_n470_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n470_), .A2(G78gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT110), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n714_), .B2(new_n735_), .ZN(G1335gat));
  AND3_X1   g535(.A1(new_n660_), .A2(new_n668_), .A3(new_n620_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT111), .A3(new_n570_), .A4(new_n539_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n660_), .A2(new_n668_), .A3(new_n570_), .A4(new_n620_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n539_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AND4_X1   g541(.A1(G85gat), .A2(new_n738_), .A3(new_n623_), .A4(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n713_), .A2(new_n539_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n623_), .A3(new_n678_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n483_), .B2(new_n745_), .ZN(G1336gat));
  NOR2_X1   g545(.A1(new_n468_), .A2(new_n482_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n742_), .A3(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n713_), .A2(new_n539_), .A3(new_n636_), .A4(new_n678_), .ZN(new_n749_));
  INV_X1    g548(.A(G92gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n293_), .A3(new_n742_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n479_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n744_), .A2(new_n678_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT51), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1338gat));
  NOR2_X1   g561(.A1(new_n470_), .A2(new_n480_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n744_), .A2(new_n678_), .A3(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n740_), .A2(new_n741_), .A3(new_n470_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n765_), .A2(KEYINPUT52), .A3(new_n360_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n737_), .A2(new_n570_), .A3(new_n539_), .A4(new_n653_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n764_), .C1(new_n766_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n601_), .A2(new_n570_), .A3(new_n606_), .A4(new_n619_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n539_), .A3(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT114), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n776_), .B2(new_n539_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n569_), .A2(new_n782_), .A3(new_n532_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n569_), .B2(new_n532_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n511_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n523_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n521_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n787_), .A2(new_n786_), .A3(new_n523_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n529_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT56), .B(new_n529_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n785_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n562_), .A2(new_n557_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n560_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n558_), .B(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n566_), .B(new_n800_), .C1(new_n802_), .C2(new_n799_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n567_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n536_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n626_), .B1(new_n797_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n781_), .B1(new_n807_), .B2(KEYINPUT57), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n796_), .A2(new_n532_), .A3(new_n804_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n796_), .A2(KEYINPUT58), .A3(new_n532_), .A4(new_n804_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n607_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(KEYINPUT57), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n805_), .B1(new_n796_), .B2(new_n785_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT117), .B(new_n815_), .C1(new_n816_), .C2(new_n626_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n808_), .A2(new_n813_), .A3(new_n814_), .A4(new_n817_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n779_), .A2(new_n780_), .B1(new_n818_), .B2(new_n620_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n662_), .A2(new_n623_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n775_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n620_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n778_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n778_), .A2(new_n823_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n780_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n820_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n821_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n569_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT119), .B1(new_n827_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(KEYINPUT59), .C1(new_n819_), .C2(new_n820_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n814_), .A2(new_n813_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n807_), .A2(KEYINPUT57), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n620_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(new_n831_), .A3(new_n623_), .A4(new_n662_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n569_), .A2(G113gat), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT120), .Z(new_n843_));
  AOI21_X1  g642(.A(new_n830_), .B1(new_n841_), .B2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g643(.A(new_n266_), .B1(new_n741_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n829_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n266_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n835_), .A2(new_n539_), .A3(new_n840_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n266_), .ZN(G1341gat));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n620_), .B1(new_n821_), .B2(new_n828_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(G127gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n775_), .B(new_n820_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n619_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT121), .A3(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT122), .B(G127gat), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n835_), .A2(new_n619_), .A3(new_n840_), .A4(new_n857_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n851_), .A2(new_n856_), .A3(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n829_), .B2(new_n626_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT123), .B(G134gat), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n659_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n841_), .B2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n293_), .A2(new_n470_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n623_), .A3(new_n468_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT124), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n819_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n569_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n539_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n619_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n867_), .B2(new_n626_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n659_), .A2(new_n298_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n867_), .B2(new_n876_), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n468_), .A2(new_n623_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n293_), .A3(new_n470_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n839_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n570_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(new_n400_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n219_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT62), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(KEYINPUT62), .B2(new_n884_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n819_), .A2(new_n879_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n741_), .A2(new_n220_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n839_), .A2(new_n539_), .A3(new_n880_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n887_), .A2(new_n888_), .B1(new_n889_), .B2(new_n220_), .ZN(G1349gat));
  NOR4_X1   g689(.A1(new_n881_), .A2(new_n216_), .A3(new_n403_), .A4(new_n620_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n619_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  INV_X1    g692(.A(new_n226_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n881_), .B2(new_n659_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n599_), .A2(new_n210_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n881_), .B2(new_n897_), .ZN(G1351gat));
  NAND2_X1  g697(.A1(new_n822_), .A2(new_n826_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n864_), .A3(new_n878_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n900_), .A2(new_n327_), .A3(new_n570_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n903_));
  INV_X1    g702(.A(new_n900_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904_), .B2(new_n569_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n902_), .A2(new_n903_), .A3(new_n905_), .ZN(G1352gat));
  NOR2_X1   g705(.A1(new_n900_), .A2(new_n741_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT127), .B(G204gat), .Z(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n907_), .B2(new_n910_), .ZN(G1353gat));
  NAND2_X1  g710(.A1(new_n904_), .A2(new_n619_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n912_), .B2(new_n913_), .ZN(G1354gat));
  AND3_X1   g715(.A1(new_n904_), .A2(G218gat), .A3(new_n607_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G218gat), .B1(new_n904_), .B2(new_n626_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1355gat));
endmodule


