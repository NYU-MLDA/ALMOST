//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n202_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n212_), .B(new_n213_), .C1(G85gat), .C2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  AOI21_X1  g015(.A(new_n208_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n214_), .B(new_n217_), .C1(new_n213_), .C2(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n221_));
  XOR2_X1   g020(.A(G71gat), .B(G78gat), .Z(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n219_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n210_), .A2(new_n229_), .A3(new_n218_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(KEYINPUT12), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT12), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n219_), .A2(new_n232_), .A3(new_n227_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G230gat), .A2(G233gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n228_), .A2(new_n230_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G120gat), .B(G148gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT5), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G176gat), .B(G204gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n239_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT13), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT65), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT13), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G15gat), .B(G22gat), .ZN(new_n257_));
  INV_X1    g056(.A(G1gat), .ZN(new_n258_));
  INV_X1    g057(.A(G8gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT14), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G1gat), .B(G8gat), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G29gat), .B(G36gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n268_), .A2(KEYINPUT66), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(KEYINPUT66), .ZN(new_n270_));
  XOR2_X1   g069(.A(G43gat), .B(G50gat), .Z(new_n271_));
  OR3_X1    g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n267_), .A2(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n256_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n267_), .A2(new_n274_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT71), .A3(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT15), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n274_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n267_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G113gat), .B(G141gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT72), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G169gat), .B(G197gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n277_), .B(new_n283_), .C1(new_n286_), .C2(new_n267_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n282_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT73), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n255_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G228gat), .ZN(new_n301_));
  INV_X1    g100(.A(G233gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n304_), .A2(KEYINPUT84), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308_));
  OAI22_X1  g107(.A1(new_n304_), .A2(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT84), .B1(new_n304_), .B2(new_n305_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n306_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n308_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT85), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n318_), .B(KEYINPUT1), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n317_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n304_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n323_), .A2(new_n307_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n314_), .A2(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT87), .B1(new_n331_), .B2(G197gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(G204gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n332_), .B(new_n335_), .C1(new_n334_), .C2(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n330_), .A2(new_n336_), .A3(KEYINPUT88), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n336_), .A2(KEYINPUT21), .ZN(new_n341_));
  INV_X1    g140(.A(new_n328_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G197gat), .B(G204gat), .Z(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(KEYINPUT21), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n339_), .A2(new_n340_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n303_), .B1(new_n327_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n340_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI221_X1 g148(.A(new_n349_), .B1(new_n301_), .B2(new_n302_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(KEYINPUT89), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n314_), .A2(new_n320_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n322_), .A2(new_n323_), .A3(new_n307_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n361_), .B2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n325_), .A2(new_n326_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G22gat), .B(G50gat), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n365_), .B(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n356_), .B1(new_n357_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n365_), .B(new_n366_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n353_), .A3(new_n371_), .A4(new_n355_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G71gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G99gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT80), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n376_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G183gat), .ZN(new_n380_));
  INV_X1    g179(.A(G190gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT23), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n380_), .A2(KEYINPUT23), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n383_), .A2(new_n386_), .A3(G183gat), .A4(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n382_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT26), .B1(new_n398_), .B2(new_n381_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT26), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G190gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n399_), .C1(new_n398_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT75), .ZN(new_n403_));
  INV_X1    g202(.A(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n407_), .A4(new_n392_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n386_), .B1(G183gat), .B2(G190gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n386_), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT76), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n412_), .B2(new_n387_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT24), .B1(new_n406_), .B2(new_n392_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT77), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n396_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT79), .B(G176gat), .Z(new_n417_));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n404_), .B2(KEYINPUT22), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT22), .B(G169gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n417_), .B(new_n419_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n382_), .A2(new_n411_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n407_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n416_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT30), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n428_), .A2(KEYINPUT81), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(KEYINPUT81), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n379_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n379_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n435_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G113gat), .B(G120gat), .Z(new_n438_));
  OR3_X1    g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT31), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n431_), .A2(new_n433_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n379_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n430_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n428_), .A2(KEYINPUT81), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n448_), .B2(new_n432_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n361_), .A2(new_n441_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n359_), .A2(new_n360_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(KEYINPUT4), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n361_), .A2(new_n454_), .A3(new_n441_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT95), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G85gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n450_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n456_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n463_), .B1(new_n456_), .B2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n444_), .A2(new_n449_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT100), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n427_), .A2(new_n349_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n380_), .A2(KEYINPUT25), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G183gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n381_), .A2(KEYINPUT26), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n401_), .A2(new_n472_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n395_), .A2(new_n408_), .A3(new_n422_), .A4(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT26), .B(G190gat), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n397_), .A2(new_n480_), .B1(new_n382_), .B2(new_n411_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n481_), .A2(KEYINPUT91), .A3(new_n395_), .A4(new_n408_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n417_), .A2(new_n420_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n407_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT92), .B1(new_n389_), .B2(new_n424_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n413_), .A2(new_n488_), .A3(new_n423_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n490_), .A3(new_n345_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT19), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n471_), .A2(new_n491_), .A3(KEYINPUT20), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT93), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT18), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G64gat), .B(G92gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NAND3_X1  g299(.A1(new_n389_), .A2(KEYINPUT92), .A3(new_n424_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n488_), .B1(new_n413_), .B2(new_n423_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n485_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n479_), .A2(new_n482_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n349_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n345_), .A2(new_n416_), .A3(new_n426_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT20), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n493_), .B(KEYINPUT90), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n427_), .B2(new_n349_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n494_), .A4(new_n491_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n496_), .A2(new_n500_), .A3(new_n510_), .A4(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n515_), .A2(KEYINPUT27), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n490_), .A2(new_n517_), .A3(new_n477_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n477_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT96), .B1(new_n503_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n520_), .A3(new_n345_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n512_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n493_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n505_), .A2(KEYINPUT20), .A3(new_n506_), .A4(new_n508_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT97), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT97), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n500_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n522_), .A2(new_n493_), .B1(KEYINPUT97), .B2(new_n524_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n500_), .B1(new_n532_), .B2(new_n525_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n515_), .A2(KEYINPUT27), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT99), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n496_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n528_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT27), .B1(new_n538_), .B2(new_n515_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n470_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  AOI211_X1 g340(.A(KEYINPUT100), .B(new_n539_), .C1(new_n531_), .C2(new_n535_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n373_), .B(new_n469_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n444_), .A2(new_n449_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n453_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n451_), .A2(new_n464_), .A3(new_n452_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n462_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT33), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n467_), .ZN(new_n549_));
  OAI211_X1 g348(.A(KEYINPUT33), .B(new_n463_), .C1(new_n456_), .C2(new_n465_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n549_), .A2(new_n538_), .A3(new_n515_), .A4(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(new_n373_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n527_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n527_), .A2(KEYINPUT98), .A3(new_n554_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n537_), .A2(new_n554_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n557_), .A2(new_n468_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n544_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n561_));
  AOI211_X1 g360(.A(new_n468_), .B(new_n539_), .C1(new_n531_), .C2(new_n535_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n373_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n543_), .A2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n300_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT36), .Z(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n286_), .A2(new_n219_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT67), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n219_), .B2(new_n274_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n274_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(new_n210_), .A3(KEYINPUT67), .A4(new_n218_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n573_), .A2(new_n570_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n569_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n229_), .B(new_n267_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT69), .B(KEYINPUT16), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n595_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n602_), .B2(new_n595_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT70), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n592_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n468_), .B(KEYINPUT101), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n565_), .A2(new_n258_), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT102), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT102), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(KEYINPUT38), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT38), .B1(new_n611_), .B2(new_n612_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n250_), .A2(new_n254_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n298_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(new_n606_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n585_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n588_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n543_), .B2(new_n563_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n258_), .B1(new_n623_), .B2(new_n468_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n613_), .A2(new_n614_), .A3(new_n624_), .ZN(G1324gat));
  AND2_X1   g424(.A1(new_n565_), .A2(new_n607_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n541_), .A2(new_n542_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n259_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n627_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(G8gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT39), .B(new_n259_), .C1(new_n623_), .C2(new_n627_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  INV_X1    g434(.A(new_n544_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G15gat), .B1(new_n622_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT41), .Z(new_n638_));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n626_), .A2(new_n639_), .A3(new_n544_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1326gat));
  NOR2_X1   g440(.A1(new_n373_), .A2(G22gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n626_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n373_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n623_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(G22gat), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n606_), .A2(new_n620_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT107), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n565_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n468_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n606_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n616_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n592_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n564_), .B2(new_n592_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n592_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n665_), .B(new_n662_), .C1(new_n543_), .C2(new_n563_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n659_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n659_), .C1(new_n664_), .C2(new_n666_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n609_), .A2(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n657_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n627_), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n627_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n300_), .A2(new_n564_), .A3(new_n654_), .A4(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT46), .B1(new_n682_), .B2(KEYINPUT108), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n674_), .B2(G36gat), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n683_), .A2(new_n687_), .ZN(G1329gat));
  NAND4_X1  g487(.A1(new_n669_), .A2(G43gat), .A3(new_n544_), .A4(new_n670_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n655_), .A2(new_n636_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(G43gat), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n656_), .B2(new_n645_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n645_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n671_), .B2(new_n694_), .ZN(G1331gat));
  AND2_X1   g494(.A1(new_n658_), .A2(new_n299_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n255_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n621_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n468_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n255_), .A2(new_n607_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT109), .Z(new_n702_));
  AOI21_X1  g501(.A(new_n298_), .B1(new_n543_), .B2(new_n563_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n608_), .A2(G57gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n700_), .B1(new_n705_), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n627_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n698_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT48), .B(new_n708_), .C1(new_n710_), .C2(new_n627_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n627_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT110), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n709_), .B(new_n717_), .C1(new_n714_), .C2(new_n711_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n698_), .B2(new_n636_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n636_), .A2(G71gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n705_), .B2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n698_), .B2(new_n373_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT50), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n373_), .A2(G78gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n705_), .B2(new_n727_), .ZN(G1335gat));
  AND2_X1   g527(.A1(new_n654_), .A2(new_n255_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n703_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n609_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n615_), .A2(new_n658_), .A3(new_n298_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n564_), .A2(new_n592_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n662_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n564_), .A2(new_n592_), .A3(new_n663_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n468_), .A2(G85gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT112), .Z(new_n740_));
  AOI21_X1  g539(.A(new_n732_), .B1(new_n738_), .B2(new_n740_), .ZN(G1336gat));
  INV_X1    g540(.A(G92gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n742_), .A3(new_n627_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(new_n627_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n742_), .ZN(G1337gat));
  NAND2_X1  g545(.A1(new_n738_), .A2(new_n544_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G99gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n544_), .A2(new_n216_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n748_), .B(new_n749_), .C1(new_n730_), .C2(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  NAND2_X1  g552(.A1(new_n736_), .A2(new_n737_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT115), .A3(new_n645_), .A4(new_n733_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(G106gat), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n645_), .B(new_n733_), .C1(new_n664_), .C2(new_n666_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n755_), .A2(new_n759_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n373_), .A2(G106gat), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OR3_X1    g562(.A1(new_n730_), .A2(KEYINPUT114), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT114), .B1(new_n730_), .B2(new_n763_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n760_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n755_), .A2(G106gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n759_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n761_), .A4(new_n766_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n768_), .A2(new_n774_), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n236_), .A2(KEYINPUT118), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n231_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n238_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT55), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n244_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n244_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT121), .B(KEYINPUT56), .C1(new_n782_), .C2(new_n244_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n281_), .A2(new_n282_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n277_), .A2(new_n282_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n293_), .B1(new_n287_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n294_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n247_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n788_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n665_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n248_), .A2(new_n793_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n783_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n784_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n298_), .B2(new_n247_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n782_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n244_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n298_), .A2(new_n805_), .A3(new_n247_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n801_), .B1(new_n804_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n620_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n800_), .B1(new_n813_), .B2(KEYINPUT120), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n799_), .B1(new_n814_), .B2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n298_), .A2(new_n805_), .A3(new_n247_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n806_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n808_), .C1(new_n803_), .C2(new_n784_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n620_), .B1(new_n819_), .B2(new_n801_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT122), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n813_), .A2(new_n800_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n606_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n826_));
  AND4_X1   g625(.A1(new_n665_), .A2(new_n696_), .A3(new_n249_), .A4(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n827_), .B(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n627_), .A2(new_n645_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n636_), .A2(new_n608_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT123), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n832_), .A2(new_n833_), .A3(new_n298_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n820_), .A2(KEYINPUT122), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n814_), .B2(new_n840_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n822_), .A2(new_n816_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n830_), .B1(new_n843_), .B2(new_n606_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT124), .B1(new_n837_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n839_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT125), .B1(new_n848_), .B2(new_n839_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n837_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n299_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n838_), .B1(new_n851_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853_));
  AOI21_X1  g652(.A(G120gat), .B1(new_n255_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n853_), .B2(G120gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n832_), .A2(new_n837_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n615_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n832_), .A2(new_n860_), .A3(new_n658_), .A4(new_n837_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n606_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n832_), .A2(new_n864_), .A3(new_n620_), .A4(new_n837_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n665_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1343gat));
  NOR4_X1   g666(.A1(new_n627_), .A2(new_n373_), .A3(new_n544_), .A4(new_n608_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n832_), .A2(new_n298_), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n832_), .A2(new_n255_), .A3(new_n868_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n832_), .A2(new_n658_), .A3(new_n868_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  NAND2_X1  g674(.A1(new_n832_), .A2(new_n868_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G162gat), .B1(new_n876_), .B2(new_n665_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n812_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n878_), .ZN(G1347gat));
  NOR4_X1   g678(.A1(new_n676_), .A2(new_n645_), .A3(new_n636_), .A4(new_n609_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n832_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n420_), .A3(new_n298_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n658_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n298_), .B(new_n880_), .C1(new_n883_), .C2(new_n830_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G169gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n832_), .A2(new_n880_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n405_), .A3(new_n615_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n881_), .A2(new_n255_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n417_), .B2(new_n892_), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n832_), .A2(new_n658_), .A3(new_n880_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n397_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n380_), .B2(new_n894_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n881_), .A2(new_n620_), .A3(new_n480_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G190gat), .B1(new_n890_), .B2(new_n665_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1351gat));
  NOR2_X1   g698(.A1(new_n544_), .A2(new_n373_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n627_), .A2(new_n699_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n832_), .A2(new_n298_), .A3(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n844_), .A2(new_n901_), .ZN(new_n905_));
  AND2_X1   g704(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n905_), .B(new_n255_), .C1(new_n906_), .C2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n832_), .A2(new_n902_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n615_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n910_), .B2(new_n907_), .ZN(G1353gat));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n905_), .B(new_n658_), .C1(new_n912_), .C2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n909_), .A2(new_n606_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n912_), .ZN(G1354gat));
  AOI211_X1 g715(.A(new_n812_), .B(new_n901_), .C1(new_n825_), .C2(new_n831_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G218gat), .B1(new_n917_), .B2(KEYINPUT127), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n909_), .B2(new_n812_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n592_), .A2(G218gat), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n918_), .A2(new_n920_), .B1(new_n905_), .B2(new_n921_), .ZN(G1355gat));
endmodule


