//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n217_), .A3(new_n213_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n218_), .A2(KEYINPUT86), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT86), .B1(new_n218_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G134gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G127gat), .ZN(new_n228_));
  INV_X1    g027(.A(G127gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G134gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n230_), .A3(KEYINPUT84), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT84), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n226_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n230_), .A3(KEYINPUT84), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n225_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n224_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT92), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n224_), .A2(new_n239_), .A3(new_n243_), .A4(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n218_), .A2(new_n221_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n218_), .A2(KEYINPUT86), .A3(new_n221_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(new_n238_), .A3(new_n233_), .A4(new_n214_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n224_), .A2(new_n239_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT4), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n246_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n246_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G57gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G8gat), .B(G36gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT19), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT80), .A4(new_n276_), .ZN(new_n280_));
  OAI21_X1  g079(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT25), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n274_), .A2(new_n276_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n285_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT21), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n285_), .A2(KEYINPUT81), .A3(new_n300_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n286_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n297_), .A2(new_n318_), .A3(new_n299_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n284_), .A2(KEYINPUT91), .A3(new_n277_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT91), .B1(new_n284_), .B2(new_n277_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n311_), .A2(new_n312_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n316_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n271_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n270_), .A2(new_n316_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n303_), .A2(new_n314_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n268_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n285_), .A2(KEYINPUT81), .A3(new_n300_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT81), .B1(new_n285_), .B2(new_n300_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n323_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n284_), .A2(new_n277_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n284_), .A2(KEYINPUT91), .A3(new_n277_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n298_), .B1(new_n286_), .B2(new_n317_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n336_), .A2(new_n337_), .B1(new_n338_), .B2(new_n297_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n313_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n270_), .B1(new_n333_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n323_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(new_n326_), .C1(new_n323_), .C2(new_n322_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n343_), .A3(new_n267_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n263_), .A2(new_n330_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n245_), .A2(new_n256_), .A3(new_n254_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n252_), .A2(new_n253_), .A3(new_n246_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n261_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n346_), .A2(KEYINPUT33), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n347_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n254_), .A2(new_n256_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n353_), .B2(new_n245_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n354_), .A2(KEYINPUT93), .A3(KEYINPUT33), .A4(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n345_), .A2(new_n351_), .A3(new_n355_), .A4(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n214_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT28), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n251_), .A2(new_n363_), .A3(new_n360_), .A4(new_n214_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G22gat), .B(G50gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n213_), .A2(new_n212_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n210_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n209_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(new_n203_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n361_), .A2(KEYINPUT28), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT87), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n368_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT90), .B1(new_n370_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT89), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(G228gat), .A3(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n386_), .B(new_n388_), .Z(new_n389_));
  AOI21_X1  g188(.A(new_n313_), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(G228gat), .B2(G233gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n323_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n386_), .B(new_n388_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n369_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n381_), .A2(new_n368_), .A3(new_n382_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n384_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n399_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n397_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT90), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n341_), .A2(new_n343_), .A3(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n333_), .A2(new_n340_), .A3(new_n270_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n319_), .A2(new_n334_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n313_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n271_), .B1(new_n342_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n348_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n416_));
  OAI221_X1 g215(.A(new_n408_), .B1(new_n414_), .B2(new_n407_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n359_), .A2(new_n406_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(G15gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G71gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT82), .B(G43gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G99gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n423_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n303_), .A2(KEYINPUT30), .A3(new_n314_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT83), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT83), .B1(new_n429_), .B2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n239_), .B(KEYINPUT31), .Z(new_n435_));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n431_), .A2(new_n426_), .B1(new_n436_), .B2(new_n435_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n434_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI211_X1 g240(.A(new_n400_), .B(new_n397_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n404_), .B1(new_n403_), .B2(KEYINPUT90), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n401_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n325_), .A2(new_n329_), .A3(new_n268_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n267_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n416_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n268_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n344_), .A3(KEYINPUT27), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(new_n356_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n444_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n418_), .A2(new_n441_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT95), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n418_), .A2(new_n453_), .A3(new_n456_), .A4(new_n441_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n448_), .A2(new_n451_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n444_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n415_), .A2(new_n416_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n441_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n455_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G190gat), .B(G218gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G134gat), .B(G162gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT36), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT72), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(KEYINPUT72), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n472_), .A2(KEYINPUT72), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n473_), .A3(new_n470_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(KEYINPUT15), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT15), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT9), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT65), .B(G92gat), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G85gat), .B(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT6), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n486_), .B1(new_n505_), .B2(new_n497_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n496_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n504_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT8), .B1(new_n512_), .B2(new_n486_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n488_), .A2(new_n495_), .A3(KEYINPUT66), .A4(new_n497_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n500_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n481_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n498_), .A2(new_n499_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n476_), .A2(new_n478_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n515_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n517_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n523_), .A2(new_n524_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT71), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n481_), .A2(new_n516_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n528_), .B1(new_n531_), .B2(new_n520_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n469_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT75), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n529_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n528_), .A3(new_n520_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n468_), .B(KEYINPUT36), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n536_), .A4(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT99), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n465_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT100), .ZN(new_n545_));
  XOR2_X1   g344(.A(G120gat), .B(G148gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n516_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n500_), .A2(new_n514_), .A3(new_n557_), .A4(new_n515_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n518_), .B2(new_n515_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT67), .ZN(new_n564_));
  INV_X1    g363(.A(G230gat), .ZN(new_n565_));
  INV_X1    g364(.A(G233gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n562_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(KEYINPUT12), .A3(new_n561_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n516_), .A2(new_n570_), .A3(new_n558_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n550_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(new_n563_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n562_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n550_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT69), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(KEYINPUT13), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n573_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G15gat), .B(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G8gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n519_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n478_), .A3(new_n476_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT78), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n595_), .A2(KEYINPUT78), .A3(new_n596_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(G229gat), .A3(G233gat), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n481_), .A2(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n587_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n593_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n558_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n621_), .B2(KEYINPUT77), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(KEYINPUT77), .B2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(KEYINPUT17), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT76), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n621_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n613_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT98), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n545_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n202_), .B1(new_n631_), .B2(new_n462_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n612_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n454_), .A2(KEYINPUT95), .B1(new_n460_), .B2(new_n463_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(new_n457_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n537_), .B(KEYINPUT73), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n535_), .A2(new_n536_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n535_), .A2(new_n536_), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n638_), .A2(KEYINPUT74), .B1(new_n639_), .B2(new_n469_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n638_), .A2(KEYINPUT74), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT37), .B1(new_n539_), .B2(new_n540_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n627_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n635_), .A2(new_n645_), .A3(new_n587_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT96), .Z(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n202_), .A3(new_n462_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n648_), .A2(KEYINPUT97), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT97), .B1(new_n648_), .B2(new_n649_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n632_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n649_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT101), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1324gat));
  NAND3_X1  g454(.A1(new_n647_), .A2(new_n589_), .A3(new_n459_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n631_), .A2(new_n459_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G8gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT39), .B(new_n589_), .C1(new_n631_), .C2(new_n459_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n656_), .B(new_n662_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  INV_X1    g465(.A(new_n441_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n647_), .A2(new_n420_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G15gat), .B1(new_n630_), .B2(new_n441_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n647_), .A2(new_n674_), .A3(new_n444_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G22gat), .B1(new_n630_), .B2(new_n406_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT42), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT42), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n542_), .A2(new_n627_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n587_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n635_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n462_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n627_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n613_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n644_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT43), .B(new_n688_), .C1(new_n634_), .C2(new_n457_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n465_), .B2(new_n644_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n687_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n462_), .A2(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n685_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n458_), .A2(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n635_), .A2(new_n682_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n459_), .A3(new_n695_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n699_), .B1(new_n705_), .B2(KEYINPUT46), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n705_), .B2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT103), .B(new_n703_), .C1(new_n704_), .C2(G36gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n704_), .A2(G36gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n703_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT103), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n705_), .A2(new_n708_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n715_), .A2(new_n699_), .A3(new_n707_), .A4(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n711_), .A2(new_n717_), .ZN(G1329gat));
  NAND3_X1  g517(.A1(new_n696_), .A2(G43gat), .A3(new_n667_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT105), .B(G43gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n683_), .B2(new_n441_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g522(.A1(new_n683_), .A2(G50gat), .A3(new_n406_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n696_), .A2(new_n444_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G50gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1331gat));
  NOR3_X1   g528(.A1(new_n587_), .A2(new_n612_), .A3(new_n627_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n545_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n461_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n612_), .B1(new_n634_), .B2(new_n457_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n645_), .A3(new_n681_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n461_), .A2(G57gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  OR3_X1    g535(.A1(new_n734_), .A2(G64gat), .A3(new_n458_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G64gat), .B1(new_n731_), .B2(new_n458_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n731_), .B2(new_n441_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n667_), .A2(new_n422_), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n743_), .A2(new_n744_), .B1(new_n734_), .B2(new_n745_), .ZN(G1334gat));
  OR3_X1    g545(.A1(new_n734_), .A2(G78gat), .A3(new_n406_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G78gat), .B1(new_n731_), .B2(new_n406_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT108), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT108), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n747_), .B1(new_n752_), .B2(new_n753_), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n680_), .A2(new_n587_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n733_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n462_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n689_), .A2(new_n691_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n681_), .A2(new_n633_), .A3(new_n627_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT109), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT110), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n462_), .A2(G85gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n758_), .B1(new_n763_), .B2(new_n765_), .ZN(G1336gat));
  INV_X1    g565(.A(new_n483_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n459_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n756_), .B2(new_n458_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT112), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n768_), .A2(new_n773_), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1337gat));
  NOR2_X1   g574(.A1(new_n493_), .A2(new_n494_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n756_), .A2(new_n441_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n759_), .A2(new_n667_), .A3(new_n761_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(G99gat), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1338gat));
  OAI21_X1  g580(.A(G106gat), .B1(new_n762_), .B2(new_n406_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n757_), .A2(new_n489_), .A3(new_n444_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n787_), .A3(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n612_), .A2(new_n581_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n567_), .A2(KEYINPUT115), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n795_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n578_), .B2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT55), .B(new_n797_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n550_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT55), .B1(new_n576_), .B2(new_n577_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n572_), .B2(new_n798_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n580_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n793_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n791_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n603_), .B1(new_n594_), .B2(new_n519_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n608_), .B1(new_n602_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n599_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n611_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n809_), .B1(new_n582_), .B2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT117), .B(new_n814_), .C1(new_n573_), .C2(new_n581_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n808_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n790_), .B1(new_n818_), .B2(new_n542_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n568_), .A2(new_n572_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n814_), .B1(new_n823_), .B2(new_n580_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n805_), .A2(new_n806_), .A3(new_n792_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n792_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n644_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT119), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n826_), .A2(new_n822_), .A3(new_n827_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n644_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT118), .B(new_n790_), .C1(new_n818_), .C2(new_n542_), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n818_), .A2(new_n542_), .A3(new_n790_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n821_), .A2(new_n834_), .A3(new_n835_), .A4(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n645_), .A2(new_n633_), .A3(new_n587_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n838_), .A2(new_n841_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n837_), .A2(new_n627_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n460_), .A2(new_n462_), .A3(new_n667_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n612_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n833_), .A2(new_n831_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n832_), .B1(new_n828_), .B2(new_n644_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n819_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n836_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n834_), .B2(new_n819_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n627_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n843_), .A2(new_n842_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n846_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n837_), .A2(new_n627_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n856_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n845_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(KEYINPUT59), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n633_), .B(new_n859_), .C1(new_n861_), .C2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n848_), .B1(new_n868_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n846_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n870_), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n587_), .B(new_n859_), .C1(new_n861_), .C2(new_n867_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n870_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n846_), .B2(new_n686_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n861_), .A2(new_n867_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n627_), .A2(KEYINPUT122), .ZN(new_n877_));
  MUX2_X1   g676(.A(KEYINPUT122), .B(new_n877_), .S(G127gat), .Z(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n876_), .B2(new_n878_), .ZN(G1342gat));
  OAI21_X1  g678(.A(new_n227_), .B1(new_n865_), .B2(new_n543_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT123), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n227_), .C1(new_n865_), .C2(new_n543_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n688_), .A2(new_n227_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n876_), .B2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n441_), .A2(new_n444_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT124), .Z(new_n889_));
  NAND2_X1  g688(.A1(new_n863_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n633_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n206_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n587_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n207_), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n627_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n890_), .B2(new_n688_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n543_), .A2(G162gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n890_), .B2(new_n899_), .ZN(G1347gat));
  NAND2_X1  g699(.A1(new_n459_), .A2(new_n461_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n901_), .A2(new_n444_), .A3(new_n441_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n857_), .A2(new_n612_), .A3(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT22), .B(G169gat), .Z(new_n904_));
  OR2_X1    g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n857_), .A2(KEYINPUT125), .A3(new_n612_), .A4(new_n902_), .ZN(new_n909_));
  AND4_X1   g708(.A1(new_n906_), .A2(new_n908_), .A3(G169gat), .A4(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(G169gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n903_), .B2(new_n907_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n906_), .B1(new_n912_), .B2(new_n909_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n905_), .B1(new_n910_), .B2(new_n913_), .ZN(G1348gat));
  NAND2_X1  g713(.A1(new_n857_), .A2(new_n902_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G176gat), .B1(new_n916_), .B2(new_n681_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n863_), .A2(new_n406_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n901_), .A2(new_n441_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n681_), .A2(G176gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n917_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  NOR3_X1   g723(.A1(new_n915_), .A2(new_n317_), .A3(new_n627_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n919_), .A2(new_n686_), .A3(new_n920_), .A4(new_n921_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n288_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n915_), .B2(new_n688_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n542_), .A2(new_n286_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n915_), .B2(new_n929_), .ZN(G1351gat));
  NOR3_X1   g729(.A1(new_n844_), .A2(new_n887_), .A3(new_n901_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n612_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n681_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n686_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n936_), .B2(new_n937_), .ZN(G1354gat));
  AND3_X1   g739(.A1(new_n931_), .A2(G218gat), .A3(new_n644_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n931_), .A2(new_n542_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n943_));
  AOI21_X1  g742(.A(G218gat), .B1(new_n942_), .B2(KEYINPUT127), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(G1355gat));
endmodule


