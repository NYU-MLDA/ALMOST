//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_, new_n992_, new_n993_;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT20), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT84), .B1(new_n208_), .B2(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(G197gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT87), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G211gat), .B(G218gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT21), .B1(new_n220_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n211_), .A2(G204gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n213_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n220_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n209_), .A2(new_n212_), .A3(new_n231_), .A4(new_n213_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n232_), .A2(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n230_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n225_), .A2(new_n237_), .ZN(new_n238_));
  NOR3_X1   g037(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT23), .A3(new_n250_), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n239_), .B(new_n243_), .C1(new_n247_), .C2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT89), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(KEYINPUT89), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n244_), .A2(new_n246_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT23), .B1(new_n249_), .B2(new_n250_), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(G183gat), .B2(G190gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(G169gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n207_), .B1(new_n238_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n214_), .A2(KEYINPUT85), .A3(new_n231_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n234_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n268_), .A2(new_n230_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n250_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n272_), .A2(KEYINPUT23), .B1(new_n246_), .B2(new_n244_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n263_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n242_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n239_), .B1(new_n276_), .B2(new_n240_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n255_), .A2(new_n253_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n277_), .B(new_n278_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n275_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n206_), .B1(new_n266_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n274_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n263_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n238_), .A2(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n252_), .A2(new_n257_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n269_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n205_), .A2(new_n207_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G8gat), .B(G36gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT18), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G64gat), .B(G92gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n281_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT20), .B1(new_n269_), .B2(new_n286_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n238_), .A2(new_n284_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n205_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n203_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n293_), .A3(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(KEYINPUT95), .A3(new_n293_), .A4(new_n299_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n296_), .A2(new_n297_), .A3(new_n205_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n269_), .B2(new_n286_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n206_), .B1(new_n308_), .B2(new_n285_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n294_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n304_), .A2(KEYINPUT27), .A3(new_n305_), .A4(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT28), .B(G22gat), .Z(new_n312_));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT1), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G155gat), .A3(G162gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G141gat), .B(G148gat), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT81), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT81), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  OR3_X1    g122(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n317_), .A2(new_n313_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n321_), .A2(new_n323_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT82), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n331_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n318_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n322_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n340_));
  INV_X1    g139(.A(G50gat), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n334_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n334_), .B2(new_n340_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n312_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n334_), .A2(new_n340_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G50gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n312_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n334_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n344_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(KEYINPUT88), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n269_), .B1(KEYINPUT29), .B2(new_n339_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n238_), .A2(KEYINPUT83), .B1(G228gat), .B2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n352_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n356_), .B(new_n357_), .Z(new_n360_));
  NOR3_X1   g159(.A1(new_n342_), .A2(new_n343_), .A3(new_n312_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n347_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n353_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n344_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n301_), .B(new_n311_), .C1(new_n359_), .C2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G127gat), .B(G134gat), .Z(new_n367_));
  XOR2_X1   g166(.A(G113gat), .B(G120gat), .Z(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT31), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT79), .B(G43gat), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n284_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n275_), .A2(KEYINPUT30), .A3(new_n279_), .ZN(new_n376_));
  INV_X1    g175(.A(G99gat), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n373_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n284_), .A2(new_n374_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT30), .B1(new_n275_), .B2(new_n279_), .ZN(new_n382_));
  OAI21_X1  g181(.A(G99gat), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n372_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G71gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n380_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT80), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n371_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n367_), .B(new_n368_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n332_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n339_), .A2(new_n369_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT91), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(G1gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G29gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(G29gat), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n403_), .A2(new_n404_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n404_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n407_), .A2(G29gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n402_), .A4(new_n408_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n395_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n398_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n339_), .A2(new_n369_), .A3(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n399_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n415_), .B1(new_n399_), .B2(new_n420_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n380_), .A2(new_n385_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n389_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(KEYINPUT80), .A3(new_n390_), .A4(new_n370_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n393_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n202_), .B1(new_n366_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n393_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n311_), .A2(new_n301_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n358_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n363_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(KEYINPUT96), .A3(new_n432_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n293_), .A2(KEYINPUT32), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n298_), .A2(new_n437_), .A3(new_n299_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(new_n423_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n399_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT93), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n294_), .B1(new_n281_), .B2(new_n289_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n397_), .A2(new_n417_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n416_), .A2(new_n398_), .A3(new_n419_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n411_), .A2(new_n414_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n302_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n444_), .B1(new_n443_), .B2(KEYINPUT93), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n442_), .B1(new_n445_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n359_), .A2(new_n365_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n433_), .A2(new_n434_), .A3(new_n423_), .ZN(new_n456_));
  OAI22_X1  g255(.A1(new_n454_), .A2(new_n455_), .B1(new_n431_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n393_), .A2(new_n427_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n429_), .A2(new_n436_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G232gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT34), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n377_), .A3(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT6), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT65), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT65), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G85gat), .ZN(new_n477_));
  INV_X1    g276(.A(G92gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT8), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n467_), .A2(new_n468_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n471_), .A2(new_n473_), .A3(new_n484_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n483_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n474_), .A2(new_n475_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n479_), .A2(KEYINPUT9), .A3(new_n480_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n480_), .A2(KEYINPUT9), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT64), .B(G106gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT10), .B(G99gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n493_), .B(new_n495_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT69), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n471_), .A2(new_n473_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT65), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT64), .B(G106gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n494_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .A4(new_n493_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n491_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n493_), .A3(new_n508_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n491_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n462_), .A2(new_n463_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n464_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n514_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n464_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n518_), .A4(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT36), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n527_), .A2(KEYINPUT36), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(KEYINPUT72), .A3(new_n528_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT98), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n459_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G230gat), .ZN(new_n539_));
  INV_X1    g338(.A(G233gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n500_), .A2(KEYINPUT66), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n488_), .A3(new_n469_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n481_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n490_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n482_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n504_), .B2(new_n469_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n548_), .B(new_n516_), .C1(new_n552_), .C2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT67), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n491_), .A2(new_n557_), .A3(new_n548_), .A4(new_n516_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT68), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n516_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n548_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n558_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT68), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n541_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n545_), .B(KEYINPUT12), .C1(new_n546_), .C2(new_n547_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n568_), .A2(new_n563_), .B1(new_n510_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n541_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n555_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G120gat), .B(G148gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G176gat), .B(G204gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n567_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(KEYINPUT71), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n567_), .B2(new_n575_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT13), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n581_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G8gat), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G22gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n387_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G15gat), .A2(G22gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G1gat), .A2(G8gat), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n596_), .A2(new_n597_), .B1(KEYINPUT14), .B2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n594_), .A2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n513_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n594_), .B(new_n599_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n514_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT75), .ZN(new_n611_));
  INV_X1    g410(.A(new_n608_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n602_), .A2(new_n513_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n513_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n604_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT76), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  AND3_X1   g420(.A1(new_n617_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n548_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(new_n602_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT16), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n628_), .A2(new_n634_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n591_), .A2(new_n625_), .A3(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n538_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n423_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G1gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n459_), .A2(new_n625_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n531_), .A2(new_n533_), .A3(new_n534_), .A4(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n529_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n524_), .A2(new_n532_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT37), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n638_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n591_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n645_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT97), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n645_), .A2(new_n656_), .A3(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n643_), .A3(new_n641_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n644_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n661_), .B2(new_n660_), .ZN(G1324gat));
  NAND3_X1  g462(.A1(new_n538_), .A2(new_n431_), .A3(new_n639_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n432_), .A2(G8gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n666_), .A2(new_n667_), .B1(new_n658_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT100), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672_));
  OAI221_X1 g471(.A(new_n672_), .B1(new_n658_), .B2(new_n669_), .C1(new_n667_), .C2(new_n666_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n671_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(new_n458_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n387_), .B1(new_n640_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT41), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n659_), .A2(new_n387_), .A3(new_n678_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1326gat));
  AOI21_X1  g481(.A(new_n595_), .B1(new_n640_), .B2(new_n455_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT102), .Z(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n684_), .A2(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n435_), .A2(G22gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT103), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n687_), .A2(new_n688_), .B1(new_n658_), .B2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n638_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n591_), .A2(new_n625_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n647_), .A2(new_n650_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n429_), .A2(new_n436_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n442_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n295_), .A2(new_n300_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT93), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT33), .B1(new_n421_), .B2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n698_), .A2(new_n700_), .A3(new_n445_), .A4(new_n450_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n697_), .A2(new_n701_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n456_), .A2(new_n431_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n458_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT43), .B(new_n694_), .C1(new_n696_), .C2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n695_), .B1(new_n705_), .B2(KEYINPUT104), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n696_), .A2(new_n704_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  INV_X1    g507(.A(new_n694_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n707_), .A2(KEYINPUT104), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT44), .B(new_n693_), .C1(new_n706_), .C2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT105), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n710_), .A3(new_n695_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(KEYINPUT44), .A4(new_n693_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n693_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723_), .B2(new_n423_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n535_), .A2(new_n692_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR4_X1   g525(.A1(new_n459_), .A2(new_n625_), .A3(new_n591_), .A4(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n423_), .A2(G29gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT106), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(G1328gat));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n727_), .A2(new_n732_), .A3(new_n431_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT45), .Z(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n432_), .B(new_n721_), .C1(new_n713_), .C2(new_n719_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT46), .B(new_n735_), .C1(new_n736_), .C2(new_n732_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n721_), .A2(new_n432_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n732_), .B1(new_n720_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n678_), .A2(G43gat), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(new_n721_), .C1(new_n713_), .C2(new_n719_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n727_), .A2(new_n678_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(G43gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n748_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n743_), .C1(new_n723_), .C2(new_n745_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n723_), .B2(new_n435_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n435_), .A2(G50gat), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT108), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n727_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n590_), .A2(new_n624_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n707_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n652_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n641_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n590_), .A2(new_n624_), .A3(new_n638_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n538_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n423_), .A2(KEYINPUT109), .ZN(new_n764_));
  MUX2_X1   g563(.A(KEYINPUT109), .B(new_n764_), .S(G57gat), .Z(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n763_), .B2(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n763_), .B2(new_n431_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT48), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n767_), .A3(new_n431_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n760_), .A2(new_n772_), .A3(new_n678_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n763_), .A2(new_n678_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G71gat), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g578(.A(G78gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n763_), .B2(new_n455_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT50), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n760_), .A2(new_n780_), .A3(new_n455_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  NOR3_X1   g583(.A1(new_n590_), .A2(new_n624_), .A3(new_n692_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n717_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n423_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT111), .B1(new_n759_), .B2(new_n726_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n707_), .A2(new_n789_), .A3(new_n725_), .A4(new_n758_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n477_), .A3(new_n641_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n792_), .ZN(G1336gat));
  OAI21_X1  g592(.A(G92gat), .B1(new_n786_), .B2(new_n432_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n478_), .A3(new_n431_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  NOR2_X1   g595(.A1(new_n458_), .A2(new_n497_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n791_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT112), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(new_n800_), .A3(new_n797_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n786_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n377_), .B1(new_n803_), .B2(new_n678_), .ZN(new_n804_));
  AND2_X1   g603(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n805_));
  OR3_X1    g604(.A1(new_n802_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n802_), .C2(new_n804_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n435_), .A2(new_n496_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n791_), .A2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT114), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n717_), .A2(new_n455_), .A3(new_n785_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G106gat), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n811_), .A2(new_n815_), .A3(new_n819_), .A4(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n550_), .A2(new_n551_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n823_), .A2(KEYINPUT8), .B1(new_n476_), .B2(new_n482_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n499_), .A2(new_n509_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n570_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n548_), .B1(new_n491_), .B2(new_n516_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(KEYINPUT12), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n822_), .B1(new_n828_), .B2(new_n573_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n563_), .A2(new_n568_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n574_), .A2(new_n830_), .A3(KEYINPUT55), .A4(new_n826_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n559_), .A2(new_n571_), .A3(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n830_), .A2(new_n556_), .A3(new_n558_), .A4(new_n826_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n572_), .B1(new_n835_), .B2(KEYINPUT116), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n832_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n584_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n621_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n606_), .A2(new_n608_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n613_), .A2(new_n615_), .A3(new_n612_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n617_), .B2(new_n839_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n829_), .A2(new_n831_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n828_), .B2(new_n564_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(new_n846_), .A3(new_n541_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n583_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n838_), .A2(new_n581_), .A3(new_n844_), .A4(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT118), .B1(new_n853_), .B2(new_n694_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n584_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n581_), .B1(new_n855_), .B2(new_n849_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT56), .B(new_n584_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n852_), .A4(new_n843_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n694_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n854_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT57), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n838_), .A2(new_n624_), .A3(new_n581_), .A4(new_n850_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n844_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n865_), .B1(new_n868_), .B2(new_n535_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n535_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n870_), .B(new_n864_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n862_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n638_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n590_), .A2(new_n651_), .A3(new_n625_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT54), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n590_), .A2(new_n651_), .A3(new_n877_), .A4(new_n625_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(KEYINPUT115), .B2(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(KEYINPUT115), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n874_), .A2(new_n882_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n366_), .A2(new_n423_), .A3(new_n458_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n624_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(KEYINPUT59), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n874_), .A2(KEYINPUT119), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n692_), .B1(new_n862_), .B2(new_n872_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n881_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n884_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n888_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G113gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n624_), .A2(KEYINPUT120), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(G113gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n887_), .B1(new_n897_), .B2(new_n901_), .ZN(G1340gat));
  OAI21_X1  g701(.A(G120gat), .B1(new_n896_), .B2(new_n590_), .ZN(new_n903_));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n886_), .B(new_n905_), .C1(KEYINPUT60), .C2(new_n904_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1341gat));
  OAI21_X1  g706(.A(G127gat), .B1(new_n896_), .B2(new_n638_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n885_), .A2(G127gat), .A3(new_n638_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1342gat));
  OAI21_X1  g709(.A(G134gat), .B1(new_n896_), .B2(new_n694_), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n885_), .A2(G134gat), .A3(new_n536_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1343gat));
  NOR4_X1   g712(.A1(new_n678_), .A2(new_n435_), .A3(new_n423_), .A4(new_n431_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n883_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n624_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n591_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n916_), .A2(new_n921_), .A3(new_n692_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n915_), .B2(new_n638_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n922_), .A2(new_n923_), .A3(new_n925_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1346gat));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n930_), .B1(new_n915_), .B2(new_n536_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n932_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n694_), .A2(new_n930_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n916_), .B2(new_n935_), .ZN(G1347gat));
  AOI21_X1  g735(.A(new_n891_), .B1(new_n873_), .B2(new_n638_), .ZN(new_n937_));
  AOI211_X1 g736(.A(KEYINPUT119), .B(new_n692_), .C1(new_n862_), .C2(new_n872_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n882_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT22), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n432_), .A2(new_n428_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n455_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n939_), .A2(new_n940_), .A3(new_n624_), .A4(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(G169gat), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n944_), .A2(KEYINPUT62), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(KEYINPUT62), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n939_), .A2(new_n948_), .A3(new_n624_), .A4(new_n943_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n949_), .A2(G169gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n946_), .B1(new_n947_), .B2(new_n950_), .ZN(G1348gat));
  INV_X1    g750(.A(new_n943_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n893_), .A2(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G176gat), .B1(new_n953_), .B2(new_n591_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n890_), .A2(new_n881_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT123), .B1(new_n955_), .B2(new_n455_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957_));
  OAI211_X1 g756(.A(new_n957_), .B(new_n435_), .C1(new_n890_), .C2(new_n881_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n958_), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n591_), .A2(G176gat), .A3(new_n941_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n954_), .B1(new_n959_), .B2(new_n960_), .ZN(G1349gat));
  NAND2_X1  g760(.A1(new_n941_), .A2(new_n692_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n956_), .B2(new_n958_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964_));
  OR2_X1    g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(G183gat), .B1(new_n963_), .B2(new_n964_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n638_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n967_));
  AOI22_X1  g766(.A1(new_n965_), .A2(new_n966_), .B1(new_n953_), .B2(new_n967_), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n953_), .A2(new_n255_), .A3(new_n537_), .ZN(new_n969_));
  INV_X1    g768(.A(G190gat), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n893_), .A2(new_n694_), .A3(new_n952_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n969_), .B1(new_n970_), .B2(new_n971_), .ZN(G1351gat));
  INV_X1    g771(.A(new_n456_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n678_), .A2(new_n432_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n883_), .A2(KEYINPUT125), .A3(new_n973_), .A4(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n973_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n955_), .B2(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n975_), .A2(new_n978_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(new_n624_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(KEYINPUT126), .B(G197gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n980_), .B(new_n981_), .ZN(G1352gat));
  NAND2_X1  g781(.A1(new_n979_), .A2(new_n591_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  NAND2_X1  g784(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n986_));
  AND4_X1   g785(.A1(new_n692_), .A2(new_n979_), .A3(new_n985_), .A4(new_n986_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n985_), .B1(new_n979_), .B2(new_n692_), .ZN(new_n988_));
  NOR2_X1   g787(.A1(new_n987_), .A2(new_n988_), .ZN(G1354gat));
  INV_X1    g788(.A(new_n979_), .ZN(new_n990_));
  OAI21_X1  g789(.A(G218gat), .B1(new_n990_), .B2(new_n694_), .ZN(new_n991_));
  INV_X1    g790(.A(G218gat), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n979_), .A2(new_n992_), .A3(new_n537_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n993_), .ZN(G1355gat));
endmodule


