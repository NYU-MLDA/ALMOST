//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n212_), .B(new_n215_), .Z(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n210_), .A2(new_n215_), .A3(new_n211_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G141gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT79), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  OR2_X1    g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OR3_X1    g038(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n244_), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT6), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(KEYINPUT6), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT68), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n242_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G85gat), .B(G92gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT8), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n241_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(new_n250_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n253_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT8), .ZN(new_n261_));
  OAI22_X1  g060(.A1(new_n252_), .A2(new_n255_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G92gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n253_), .B1(KEYINPUT9), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G85gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(KEYINPUT67), .A2(G92gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT67), .A2(G92gat), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT66), .B(KEYINPUT9), .Z(new_n269_));
  OAI21_X1  g068(.A(new_n264_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT65), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274_));
  AND2_X1   g073(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G106gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n248_), .A2(new_n251_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n239_), .B1(new_n262_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT12), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT68), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT68), .B1(new_n249_), .B2(new_n250_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n258_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n254_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n253_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n259_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n242_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT8), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n279_), .A2(new_n278_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n290_), .A2(new_n294_), .B1(new_n295_), .B2(new_n270_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT69), .B(new_n286_), .C1(new_n296_), .C2(new_n239_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT64), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n239_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n285_), .A2(new_n297_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n303_), .B2(new_n283_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G120gat), .B(G148gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G176gat), .B(G204gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n305_), .A2(new_n310_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT13), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n305_), .A2(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n311_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT71), .B1(new_n315_), .B2(new_n319_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n330_));
  OR3_X1    g129(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT81), .ZN(new_n335_));
  AOI211_X1 g134(.A(new_n333_), .B(new_n335_), .C1(G169gat), .C2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n333_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  INV_X1    g138(.A(G190gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT26), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G190gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n338_), .B(new_n341_), .C1(new_n342_), .C2(new_n339_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n327_), .B(KEYINPUT23), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n332_), .B1(new_n336_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT82), .B(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n346_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G134gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT83), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G113gat), .B(G120gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n351_), .A2(KEYINPUT83), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(KEYINPUT83), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(KEYINPUT84), .A3(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n350_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(G15gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT30), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT31), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n350_), .A2(new_n362_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n363_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(G78gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(new_n279_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G22gat), .B(G50gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G155gat), .B(G162gat), .Z(new_n381_));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G141gat), .A2(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT2), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n381_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n389_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(KEYINPUT29), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT28), .ZN(new_n400_));
  XOR2_X1   g199(.A(G211gat), .B(G218gat), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT21), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(KEYINPUT86), .ZN(new_n408_));
  INV_X1    g207(.A(G204gat), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n409_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(KEYINPUT21), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n406_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n398_), .A2(KEYINPUT29), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n400_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n400_), .A2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n380_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n419_), .A3(new_n379_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n362_), .A2(new_n398_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT92), .Z(new_n430_));
  AOI22_X1  g229(.A1(new_n360_), .A2(new_n361_), .B1(new_n389_), .B2(new_n397_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n398_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n428_), .B(new_n430_), .C1(new_n433_), .C2(new_n427_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n430_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n441_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT93), .B1(new_n447_), .B2(KEYINPUT33), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n428_), .B1(new_n433_), .B2(new_n427_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n435_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n441_), .B1(new_n433_), .B2(new_n430_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n447_), .A2(KEYINPUT33), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT19), .ZN(new_n456_));
  INV_X1    g255(.A(new_n332_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n335_), .B1(G169gat), .B2(G176gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n458_), .A2(new_n460_), .B1(new_n342_), .B2(new_n338_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n334_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n344_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT89), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n465_), .A3(new_n344_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n457_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n407_), .A2(new_n411_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT87), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n405_), .B1(new_n470_), .B2(new_n413_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT20), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n416_), .A2(new_n346_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n456_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G8gat), .B(G36gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n456_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n416_), .A2(new_n346_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n474_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n479_), .B1(new_n474_), .B2(new_n484_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n454_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n474_), .A2(new_n484_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n479_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(KEYINPUT91), .A3(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n449_), .A2(new_n453_), .A3(new_n487_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n474_), .A2(new_n494_), .A3(new_n484_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n472_), .A2(new_n473_), .A3(new_n456_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n482_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n434_), .A2(new_n436_), .A3(new_n446_), .ZN(new_n499_));
  OAI221_X1 g298(.A(new_n495_), .B1(new_n498_), .B2(new_n494_), .C1(new_n499_), .C2(new_n447_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n425_), .B1(new_n493_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n499_), .B2(new_n447_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n434_), .A2(new_n436_), .A3(new_n446_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n442_), .A2(KEYINPUT94), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT27), .B(new_n491_), .C1(new_n498_), .C2(new_n479_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n422_), .A2(new_n424_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n506_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n373_), .B1(new_n501_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n425_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n506_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT95), .A4(new_n372_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n372_), .A2(new_n505_), .A3(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  AOI211_X1 g320(.A(new_n232_), .B(new_n324_), .C1(new_n513_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n262_), .A2(new_n282_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n220_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT73), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n296_), .A2(new_n215_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G190gat), .B(G218gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT74), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT36), .Z(new_n539_));
  NAND4_X1  g338(.A1(new_n525_), .A2(new_n524_), .A3(new_n529_), .A4(new_n531_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n534_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n541_), .A2(new_n544_), .A3(KEYINPUT37), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n539_), .B(KEYINPUT76), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n534_), .A3(new_n540_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n548_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n545_), .B1(new_n551_), .B2(KEYINPUT37), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n212_), .B(new_n239_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT16), .ZN(new_n557_));
  XOR2_X1   g356(.A(G183gat), .B(G211gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n555_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n561_), .B2(new_n555_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT78), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n552_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n522_), .A2(new_n203_), .A3(new_n506_), .A4(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT38), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT96), .B1(new_n324_), .B2(new_n232_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n320_), .B(new_n321_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n231_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n571_), .A2(new_n574_), .A3(new_n565_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n541_), .A2(new_n544_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT97), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n515_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n568_), .A2(new_n569_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n570_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT98), .ZN(G1324gat));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n579_), .A3(new_n510_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G8gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT39), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n522_), .A2(new_n567_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n204_), .A3(new_n510_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(G1325gat));
  OAI21_X1  g392(.A(G15gat), .B1(new_n580_), .B2(new_n373_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT101), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n589_), .A2(new_n365_), .A3(new_n372_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n597_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(G1326gat));
  OR3_X1    g400(.A1(new_n588_), .A2(G22gat), .A3(new_n511_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n575_), .A2(new_n425_), .A3(new_n579_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT42), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(G22gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n603_), .B2(G22gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(G1327gat));
  NOR2_X1   g406(.A1(new_n577_), .A2(new_n565_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n522_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n506_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n571_), .A2(new_n574_), .A3(new_n566_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n552_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n552_), .B2(new_n615_), .ZN(new_n616_));
  AOI211_X1 g415(.A(new_n613_), .B(new_n616_), .C1(new_n513_), .C2(new_n521_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n445_), .A2(new_n448_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n453_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n500_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n512_), .B1(new_n621_), .B2(new_n511_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n521_), .B1(new_n622_), .B2(new_n372_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n618_), .B1(new_n623_), .B2(new_n552_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n612_), .B(KEYINPUT44), .C1(new_n617_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT44), .B1(new_n627_), .B2(KEYINPUT103), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n612_), .B(new_n629_), .C1(new_n617_), .C2(new_n624_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n626_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n506_), .A2(G29gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n611_), .B1(new_n631_), .B2(new_n632_), .ZN(G1328gat));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(G36gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n631_), .B2(new_n510_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n610_), .A2(new_n636_), .A3(new_n510_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT45), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n571_), .A2(new_n574_), .A3(new_n566_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n623_), .A2(new_n552_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n616_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n623_), .A2(new_n552_), .A3(new_n618_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n647_), .B2(new_n629_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n630_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n510_), .B(new_n625_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n635_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n641_), .A2(new_n654_), .ZN(G1329gat));
  INV_X1    g454(.A(G43gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n373_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n631_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n609_), .B2(new_n373_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT47), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1330gat));
  OR3_X1    g463(.A1(new_n609_), .A2(G50gat), .A3(new_n511_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n631_), .A2(new_n666_), .A3(new_n425_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G50gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n631_), .B2(new_n425_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1331gat));
  AOI21_X1  g469(.A(new_n231_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT106), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n324_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n567_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G57gat), .B1(new_n675_), .B2(new_n506_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n572_), .A2(new_n566_), .A3(new_n231_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n579_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(G57gat), .A3(new_n506_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT107), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1332gat));
  INV_X1    g480(.A(G64gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n678_), .B2(new_n510_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT48), .Z(new_n684_));
  NAND2_X1  g483(.A1(new_n510_), .A2(new_n682_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n674_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n678_), .B2(new_n372_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n372_), .A2(new_n687_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n674_), .B2(new_n690_), .ZN(G1334gat));
  NAND2_X1  g490(.A1(new_n678_), .A2(new_n425_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G78gat), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT50), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(KEYINPUT50), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n425_), .A2(new_n375_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT109), .Z(new_n701_));
  OAI211_X1 g500(.A(new_n698_), .B(new_n699_), .C1(new_n674_), .C2(new_n701_), .ZN(G1335gat));
  NAND2_X1  g501(.A1(new_n673_), .A2(new_n608_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n265_), .A3(new_n506_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n565_), .A2(new_n231_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n324_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT110), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n324_), .A2(new_n709_), .A3(new_n706_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n645_), .A2(new_n646_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n506_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n705_), .B1(new_n265_), .B2(new_n713_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n704_), .B2(new_n510_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n266_), .A2(new_n267_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n510_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n711_), .B2(new_n718_), .ZN(G1337gat));
  NAND2_X1  g518(.A1(new_n711_), .A2(new_n372_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G99gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n372_), .A2(new_n278_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n703_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g523(.A1(new_n673_), .A2(new_n279_), .A3(new_n425_), .A4(new_n608_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n708_), .A2(new_n710_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n425_), .B(new_n727_), .C1(new_n617_), .C2(new_n624_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n728_), .B2(G106gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n726_), .A3(G106gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n726_), .B(new_n733_), .C1(new_n728_), .C2(G106gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n725_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n725_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  NAND3_X1  g538(.A1(new_n285_), .A2(new_n301_), .A3(new_n297_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n299_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT55), .A3(new_n302_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n285_), .A2(new_n301_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n300_), .A4(new_n297_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n742_), .A2(new_n743_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n743_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT56), .B(new_n310_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n742_), .A2(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n742_), .A2(new_n743_), .A3(new_n746_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(KEYINPUT56), .A4(new_n310_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n310_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n216_), .A2(new_n217_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n221_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n228_), .A3(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT115), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT115), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n229_), .A3(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n313_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n767_), .A3(KEYINPUT58), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n552_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n231_), .A2(new_n316_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n759_), .B2(new_n749_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n766_), .A2(new_n314_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n577_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT57), .B(new_n577_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n566_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n566_), .A2(new_n231_), .A3(new_n320_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n613_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT54), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n514_), .A2(new_n506_), .A3(new_n372_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT117), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G113gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n231_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n232_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(new_n790_), .ZN(G1340gat));
  AOI21_X1  g595(.A(new_n572_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n797_));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n800_));
  AOI21_X1  g599(.A(G120gat), .B1(new_n324_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n800_), .B2(G120gat), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n789_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n799_), .B1(new_n789_), .B2(new_n802_), .ZN(new_n804_));
  OAI22_X1  g603(.A1(new_n797_), .A2(new_n798_), .B1(new_n803_), .B2(new_n804_), .ZN(G1341gat));
  INV_X1    g604(.A(G127gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n789_), .A2(new_n806_), .A3(new_n565_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n566_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n806_), .ZN(G1342gat));
  AOI21_X1  g608(.A(G134gat), .B1(new_n789_), .B2(new_n578_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n792_), .A2(new_n794_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n552_), .A2(G134gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT119), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n811_), .B2(new_n813_), .ZN(G1343gat));
  NOR2_X1   g613(.A1(new_n511_), .A2(new_n372_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n506_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n232_), .ZN(new_n819_));
  INV_X1    g618(.A(G141gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1344gat));
  NOR2_X1   g620(.A1(new_n818_), .A2(new_n572_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT120), .B(G148gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  NOR2_X1   g623(.A1(new_n818_), .A2(new_n566_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n825_), .B(new_n827_), .ZN(G1346gat));
  OAI21_X1  g627(.A(G162gat), .B1(new_n818_), .B2(new_n613_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n577_), .A2(G162gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n818_), .B2(new_n830_), .ZN(G1347gat));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n832_));
  INV_X1    g631(.A(G169gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n372_), .A3(new_n231_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT121), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n425_), .B(new_n836_), .C1(new_n781_), .C2(new_n784_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n833_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n836_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n773_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n310_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n749_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n775_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n846_), .B2(new_n577_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n779_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n770_), .A2(new_n552_), .A3(new_n771_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n565_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n783_), .B(KEYINPUT54), .Z(new_n852_));
  OAI211_X1 g651(.A(new_n511_), .B(new_n840_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n832_), .B1(new_n839_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G169gat), .B1(new_n853_), .B2(KEYINPUT122), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n425_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n838_), .B1(new_n857_), .B2(new_n840_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n858_), .A3(KEYINPUT62), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n372_), .A3(new_n834_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT22), .B(G169gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n231_), .A2(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT123), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n855_), .A2(new_n859_), .B1(new_n860_), .B2(new_n863_), .ZN(G1348gat));
  NOR2_X1   g663(.A1(new_n860_), .A2(new_n572_), .ZN(new_n865_));
  INV_X1    g664(.A(G176gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1349gat));
  INV_X1    g666(.A(new_n860_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G183gat), .B1(new_n868_), .B2(new_n565_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n860_), .A2(new_n338_), .A3(new_n566_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n860_), .B2(new_n613_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n578_), .A2(new_n342_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n860_), .B2(new_n873_), .ZN(G1351gat));
  OAI211_X1 g673(.A(new_n815_), .B(new_n834_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n231_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g677(.A1(new_n817_), .A2(new_n409_), .A3(new_n324_), .A4(new_n834_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n817_), .A2(KEYINPUT124), .A3(new_n324_), .A4(new_n834_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n785_), .A2(new_n324_), .A3(new_n815_), .A4(new_n834_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n409_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n881_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n875_), .B2(new_n572_), .ZN(new_n887_));
  AND4_X1   g686(.A1(KEYINPUT125), .A2(new_n887_), .A3(G204gat), .A4(new_n882_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n566_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT126), .B1(new_n875_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n817_), .A2(new_n893_), .A3(new_n834_), .A4(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI21_X1  g697(.A(G218gat), .B1(new_n875_), .B2(new_n613_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n875_), .A2(G218gat), .A3(new_n577_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n901_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(KEYINPUT127), .A3(new_n899_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1355gat));
endmodule


