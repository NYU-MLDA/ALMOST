//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT20), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT97), .ZN(new_n207_));
  INV_X1    g006(.A(G211gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(G218gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(G211gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(G211gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(G218gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT97), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT99), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT99), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT95), .ZN(new_n220_));
  INV_X1    g019(.A(G197gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(G204gat), .ZN(new_n222_));
  INV_X1    g021(.A(G204gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n222_), .A2(new_n224_), .B1(new_n221_), .B2(G204gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(new_n219_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT94), .B1(new_n223_), .B2(G197gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(new_n221_), .B2(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT94), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n221_), .A3(G204gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n223_), .A2(KEYINPUT93), .A3(G197gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n230_), .A2(new_n232_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(KEYINPUT21), .A2(new_n236_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n221_), .A2(G204gat), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n223_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT95), .B1(new_n223_), .B2(G197gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n226_), .B(new_n238_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT96), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT96), .B1(new_n225_), .B2(new_n226_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT98), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n225_), .A2(KEYINPUT96), .A3(new_n226_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT98), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n237_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n229_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT85), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G183gat), .A3(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT23), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G183gat), .A3(G190gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT100), .B(KEYINPUT24), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n257_), .A2(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT101), .ZN(new_n263_));
  AND2_X1   g062(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G190gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT26), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(KEYINPUT26), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n261_), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(new_n260_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n262_), .B2(KEYINPUT101), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n272_), .A2(KEYINPUT22), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(KEYINPUT22), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n273_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n274_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT102), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n253_), .A2(new_n258_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n254_), .A2(new_n256_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n258_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n263_), .A2(new_n278_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n206_), .B1(new_n252_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n272_), .A2(new_n273_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT24), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n275_), .B2(KEYINPUT24), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n269_), .A2(new_n268_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT84), .B(G183gat), .Z(new_n296_));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n298_), .B2(new_n265_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n257_), .A2(new_n259_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n267_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n279_), .A2(new_n280_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(G176gat), .B1(new_n280_), .B2(KEYINPUT86), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n274_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n294_), .A2(new_n299_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n252_), .A2(KEYINPUT103), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT103), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n249_), .A2(new_n250_), .A3(new_n237_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n250_), .B1(new_n249_), .B2(new_n237_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n228_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n308_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n205_), .B(new_n290_), .C1(new_n309_), .C2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT104), .B(KEYINPUT18), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  OAI211_X1 g120(.A(new_n308_), .B(new_n228_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(KEYINPUT20), .C1(new_n252_), .C2(new_n289_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n204_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n316_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n316_), .B2(new_n324_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n202_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT111), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT111), .B(new_n202_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n316_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT27), .ZN(new_n333_));
  INV_X1    g132(.A(new_n321_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT110), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n323_), .B2(new_n204_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n278_), .A2(new_n263_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n284_), .A2(new_n288_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n206_), .B1(new_n313_), .B2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT110), .A3(new_n205_), .A4(new_n322_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT103), .B1(new_n252_), .B2(new_n308_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n313_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n336_), .B(new_n341_), .C1(new_n345_), .C2(new_n205_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n333_), .B1(new_n334_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT91), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(G155gat), .B2(G162gat), .ZN(new_n352_));
  INV_X1    g151(.A(G141gat), .ZN(new_n353_));
  INV_X1    g152(.A(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT3), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT2), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(KEYINPUT3), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n359_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT1), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n357_), .B(new_n355_), .C1(new_n351_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT29), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n313_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G228gat), .ZN(new_n370_));
  INV_X1    g169(.A(G233gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n313_), .B(new_n368_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT92), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n367_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT28), .B1(new_n367_), .B2(KEYINPUT29), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G22gat), .B(G50gat), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n380_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n308_), .B(KEYINPUT30), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(G15gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT87), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n392_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n388_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(KEYINPUT89), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(KEYINPUT89), .ZN(new_n399_));
  XOR2_X1   g198(.A(G113gat), .B(G120gat), .Z(new_n400_));
  OR3_X1    g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT31), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT88), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n396_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n396_), .A2(new_n405_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n367_), .A2(new_n403_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n363_), .A2(new_n401_), .A3(new_n366_), .A4(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT4), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT105), .Z(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n367_), .A2(new_n403_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT106), .B(KEYINPUT0), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT107), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n420_), .B(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n408_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n331_), .A2(new_n348_), .A3(new_n387_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT112), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n347_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(KEYINPUT112), .A3(new_n387_), .A4(new_n430_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n408_), .B(KEYINPUT90), .Z(new_n436_));
  INV_X1    g235(.A(new_n380_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n386_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n429_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n316_), .A2(new_n324_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT109), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT109), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n316_), .A2(new_n444_), .A3(new_n324_), .A4(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n441_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n428_), .B1(new_n346_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n325_), .A2(new_n326_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n452_));
  INV_X1    g251(.A(new_n411_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT108), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n415_), .A2(new_n417_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n409_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n456_), .A2(new_n424_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n451_), .A2(new_n452_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n450_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n434_), .A2(new_n440_), .B1(new_n462_), .B2(new_n387_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n433_), .B(new_n435_), .C1(new_n436_), .C2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT13), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G230gat), .A2(G233gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT6), .ZN(new_n468_));
  OAI22_X1  g267(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G85gat), .B(G92gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(KEYINPUT66), .A3(new_n474_), .A4(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n488_));
  INV_X1    g287(.A(G85gat), .ZN(new_n489_));
  INV_X1    g288(.A(G92gat), .ZN(new_n490_));
  OR3_X1    g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT9), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n487_), .A2(new_n488_), .A3(new_n468_), .A4(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G78gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(KEYINPUT11), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT67), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n493_), .B(new_n497_), .C1(KEYINPUT11), .C2(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n484_), .B(new_n492_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT12), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n482_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n492_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n484_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(KEYINPUT68), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT69), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n492_), .B(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n504_), .A2(KEYINPUT12), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT70), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n513_), .B1(new_n505_), .B2(KEYINPUT68), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n509_), .B(new_n482_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n515_), .B(KEYINPUT70), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n466_), .B(new_n508_), .C1(new_n516_), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n502_), .A2(new_n507_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n466_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G120gat), .B(G148gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NAND3_X1  g328(.A1(new_n521_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n465_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT13), .A3(new_n530_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT15), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540_));
  INV_X1    g339(.A(G1gat), .ZN(new_n541_));
  INV_X1    g340(.A(G8gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT79), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n547_), .B(new_n549_), .ZN(new_n550_));
  MUX2_X1   g349(.A(new_n538_), .B(new_n539_), .S(new_n550_), .Z(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n550_), .B(new_n538_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G113gat), .B(G141gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT83), .ZN(new_n558_));
  XOR2_X1   g357(.A(G169gat), .B(G197gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n556_), .B(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n533_), .A2(new_n535_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n464_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n514_), .A2(new_n539_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n505_), .A2(new_n506_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n538_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT74), .Z(new_n574_));
  NAND4_X1  g373(.A1(new_n566_), .A2(new_n567_), .A3(new_n572_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n574_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n539_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n492_), .B(KEYINPUT69), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n484_), .B2(new_n509_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n579_), .B2(new_n511_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT75), .B1(new_n576_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n573_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n514_), .A2(new_n584_), .A3(new_n539_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n484_), .A2(new_n492_), .A3(new_n538_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT73), .B1(new_n586_), .B2(new_n570_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n572_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n580_), .A2(new_n584_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n583_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n582_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n595_), .B(KEYINPUT36), .Z(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT76), .Z(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n582_), .B2(new_n592_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT77), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT77), .B(new_n599_), .C1(new_n582_), .C2(new_n592_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n582_), .A2(new_n592_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n598_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n597_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n605_), .B1(new_n608_), .B2(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n607_), .A2(KEYINPUT78), .A3(new_n610_), .A4(new_n597_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n604_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT80), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT17), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT82), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n550_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(new_n504_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT81), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n617_), .A2(new_n618_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n612_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n565_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n541_), .A3(new_n429_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT113), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n563_), .A2(KEYINPUT114), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT114), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n533_), .A2(new_n535_), .A3(new_n638_), .A4(new_n562_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n630_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT115), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n640_), .A2(KEYINPUT115), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n464_), .A2(new_n608_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n429_), .A3(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n633_), .A2(new_n634_), .B1(G1gat), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n636_), .A2(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(new_n434_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n632_), .A2(new_n542_), .A3(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n650_), .A3(new_n646_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(G8gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n652_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT40), .B(new_n651_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(KEYINPUT116), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n645_), .A2(new_n646_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n436_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G15gat), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT41), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n632_), .A2(new_n390_), .A3(new_n436_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n665_), .B2(KEYINPUT41), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n662_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n665_), .A2(KEYINPUT41), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(KEYINPUT116), .A3(new_n666_), .A4(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1326gat));
  OAI21_X1  g472(.A(G22gat), .B1(new_n663_), .B2(new_n387_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT117), .B(KEYINPUT42), .Z(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n387_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n632_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n677_), .A3(new_n680_), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n641_), .A2(new_n608_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n565_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n429_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n640_), .A2(new_n630_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n464_), .A2(new_n688_), .A3(new_n612_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n464_), .B2(new_n612_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n687_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(G29gat), .A3(new_n429_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n464_), .A2(new_n612_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n464_), .A2(new_n688_), .A3(new_n612_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n686_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT118), .B(KEYINPUT44), .Z(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n685_), .B1(new_n692_), .B2(new_n699_), .ZN(G1328gat));
  OAI211_X1 g499(.A(new_n691_), .B(new_n650_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n434_), .A2(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n565_), .A2(new_n682_), .A3(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n408_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n691_), .B(new_n712_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n683_), .B2(new_n664_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n684_), .B2(new_n679_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n691_), .A2(G50gat), .A3(new_n679_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n699_), .ZN(G1331gat));
  NAND2_X1  g518(.A1(new_n464_), .A2(new_n608_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n533_), .A2(new_n535_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR4_X1   g521(.A1(new_n720_), .A2(new_n630_), .A3(new_n562_), .A4(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(G57gat), .A3(new_n429_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT119), .ZN(new_n725_));
  INV_X1    g524(.A(new_n562_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n464_), .A2(new_n726_), .A3(new_n721_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(new_n631_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n429_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1332gat));
  INV_X1    g529(.A(G64gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n723_), .B2(new_n650_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT48), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(new_n731_), .A3(new_n650_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n723_), .B2(new_n436_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT49), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n736_), .A3(new_n436_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n723_), .B2(new_n679_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n728_), .A2(new_n741_), .A3(new_n679_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  AND2_X1   g544(.A1(new_n727_), .A2(new_n682_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n489_), .A3(new_n429_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n694_), .A2(new_n695_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n722_), .A2(new_n641_), .A3(new_n562_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n429_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n747_), .B1(new_n753_), .B2(new_n489_), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n490_), .A3(new_n650_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n650_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n757_), .B2(new_n490_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n750_), .B2(new_n664_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n746_), .A2(new_n485_), .A3(new_n407_), .A4(new_n406_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n746_), .A2(new_n486_), .A3(new_n679_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n679_), .B(new_n749_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G106gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G106gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n763_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  NAND3_X1  g571(.A1(new_n604_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n721_), .A2(new_n630_), .A3(new_n562_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(KEYINPUT54), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT120), .B1(new_n521_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT70), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n785_), .A2(new_n519_), .B1(new_n507_), .B2(new_n503_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT55), .A4(new_n466_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n782_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT55), .B1(new_n786_), .B2(new_n466_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n786_), .A2(new_n466_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n529_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n556_), .A2(new_n561_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n555_), .A2(new_n552_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n560_), .C1(new_n552_), .C2(new_n551_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n531_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n793_), .A2(new_n794_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n780_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n789_), .A2(new_n792_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n529_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n795_), .A4(new_n800_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(new_n612_), .A3(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n799_), .B1(new_n534_), .B2(new_n530_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n562_), .A2(new_n530_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n794_), .A2(KEYINPUT121), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n793_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n521_), .A2(new_n781_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n508_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n523_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n782_), .B2(new_n788_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n813_), .B1(new_n820_), .B2(new_n529_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n811_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n608_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n810_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n811_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n804_), .A2(new_n805_), .A3(new_n814_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n812_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n793_), .A2(new_n814_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n810_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n608_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n809_), .A2(new_n824_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n779_), .B1(new_n833_), .B2(new_n630_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n650_), .A2(new_n679_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n408_), .A2(new_n428_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n562_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n837_), .B(KEYINPUT123), .Z(new_n842_));
  OR3_X1    g641(.A1(new_n834_), .A2(KEYINPUT59), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n834_), .B2(new_n838_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n843_), .A2(new_n562_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n845_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n721_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n839_), .A2(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n843_), .A2(new_n721_), .A3(new_n844_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n848_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n839_), .A2(new_n854_), .A3(new_n641_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n843_), .A2(new_n641_), .A3(new_n844_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(G1342gat));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n839_), .A2(new_n858_), .A3(new_n823_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n843_), .A2(new_n612_), .A3(new_n844_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1343gat));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n833_), .A2(new_n630_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n779_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n664_), .A2(new_n679_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(new_n650_), .A3(new_n428_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n867_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n834_), .A2(KEYINPUT124), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n562_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G141gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n865_), .A2(new_n862_), .A3(new_n867_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT124), .B1(new_n834_), .B2(new_n869_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n353_), .A3(new_n562_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n876_), .ZN(G1344gat));
  OAI21_X1  g676(.A(new_n721_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G148gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n354_), .A3(new_n721_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n875_), .B2(new_n641_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n882_), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n630_), .B(new_n884_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n875_), .A2(new_n887_), .A3(new_n823_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n773_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n664_), .A2(KEYINPUT125), .A3(new_n434_), .A4(new_n429_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n434_), .A2(new_n429_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n436_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n387_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n865_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n726_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n891_), .B1(new_n899_), .B2(new_n272_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT62), .B(G169gat), .C1(new_n898_), .C2(new_n726_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n280_), .A3(new_n279_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(new_n896_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n721_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g705(.A(new_n296_), .B1(new_n904_), .B2(new_n641_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n266_), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n834_), .A2(new_n630_), .A3(new_n908_), .A4(new_n896_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT126), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(new_n641_), .A3(new_n266_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n834_), .A2(new_n630_), .A3(new_n896_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(new_n912_), .C1(new_n913_), .C2(new_n296_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n898_), .B2(new_n773_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n904_), .A2(new_n823_), .A3(new_n295_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n866_), .A2(new_n434_), .A3(new_n429_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n865_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n726_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n221_), .ZN(G1352gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n722_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n223_), .ZN(G1353gat));
  XOR2_X1   g723(.A(KEYINPUT63), .B(G211gat), .Z(new_n925_));
  NAND4_X1  g724(.A1(new_n865_), .A2(new_n641_), .A3(new_n919_), .A4(new_n925_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n926_), .A2(KEYINPUT127), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(KEYINPUT127), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n920_), .B2(new_n630_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n920_), .B2(new_n773_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n823_), .A2(new_n210_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n920_), .B2(new_n933_), .ZN(G1355gat));
endmodule


