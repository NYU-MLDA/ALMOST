//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n988_, new_n989_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT84), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n212_), .A2(new_n213_), .A3(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n206_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(new_n210_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT84), .ZN(new_n223_));
  OAI21_X1  g022(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(new_n223_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G190gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT24), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n238_), .A2(KEYINPUT83), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT83), .B1(new_n238_), .B2(new_n239_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n208_), .A2(new_n210_), .B1(new_n242_), .B2(new_n239_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n236_), .A2(new_n240_), .A3(new_n241_), .A4(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n228_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G197gat), .B(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G211gat), .ZN(new_n250_));
  INV_X1    g049(.A(G211gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G218gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G204gat), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G197gat), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n256_), .A2(new_n258_), .A3(KEYINPUT92), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT21), .B1(new_n256_), .B2(KEYINPUT92), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n248_), .B(new_n254_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n246_), .A2(new_n247_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n253_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n245_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n227_), .B1(new_n271_), .B2(KEYINPUT98), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT98), .ZN(new_n273_));
  AOI211_X1 g072(.A(new_n273_), .B(new_n270_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n274_));
  AND2_X1   g073(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n229_), .B(new_n231_), .C1(new_n275_), .C2(new_n235_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n243_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT97), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n237_), .A2(new_n278_), .A3(KEYINPUT24), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n237_), .B2(KEYINPUT24), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n239_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n272_), .A2(new_n274_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n265_), .B(new_n269_), .C1(new_n264_), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n264_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n253_), .B1(new_n247_), .B2(new_n246_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n256_), .A2(new_n258_), .A3(KEYINPUT92), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n257_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT21), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n285_), .A2(new_n288_), .B1(new_n253_), .B2(new_n262_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n228_), .A2(new_n244_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n290_), .A3(KEYINPUT20), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n291_), .A2(KEYINPUT99), .A3(new_n267_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT99), .B1(new_n291_), .B2(new_n267_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n205_), .B(new_n283_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n267_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT99), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(KEYINPUT99), .A3(new_n267_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(KEYINPUT100), .A3(new_n205_), .A4(new_n283_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n283_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n205_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G113gat), .B(G120gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(G141gat), .ZN(new_n310_));
  INV_X1    g109(.A(G148gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G155gat), .ZN(new_n313_));
  INV_X1    g112(.A(G162gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT87), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n315_), .A2(new_n317_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n312_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n317_), .ZN(new_n328_));
  NOR4_X1   g127(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n328_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n309_), .B1(new_n327_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT3), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n331_), .A2(new_n332_), .A3(new_n330_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n324_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n307_), .B(new_n308_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n322_), .A2(new_n321_), .A3(new_n319_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n348_), .A2(new_n318_), .B1(new_n325_), .B2(new_n324_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n346_), .B(new_n347_), .C1(new_n349_), .C2(new_n312_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n350_), .A3(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n354_), .B(new_n309_), .C1(new_n327_), .C2(new_n340_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n341_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(KEYINPUT33), .A3(new_n357_), .A4(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n341_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n368_), .A2(KEYINPUT101), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT101), .B1(new_n368_), .B2(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n283_), .B(new_n373_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n291_), .A2(new_n267_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT102), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n261_), .A2(new_n377_), .A3(new_n263_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n282_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n376_), .B1(new_n380_), .B2(new_n268_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n264_), .A2(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n289_), .A2(new_n377_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT102), .B(KEYINPUT20), .C1(new_n384_), .C2(new_n282_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n265_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n375_), .B1(new_n386_), .B2(new_n267_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n374_), .B1(new_n387_), .B2(new_n373_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n356_), .A2(new_n357_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n364_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT103), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n368_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(KEYINPUT103), .A3(new_n364_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n306_), .A2(new_n372_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n323_), .A2(new_n326_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n312_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n346_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT29), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT91), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .A4(new_n384_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n264_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414_));
  INV_X1    g213(.A(G22gat), .ZN(new_n415_));
  INV_X1    g214(.A(G50gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G22gat), .A2(G50gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT28), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT28), .B1(new_n417_), .B2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT90), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  AND4_X1   g225(.A1(new_n414_), .A2(new_n398_), .A3(new_n426_), .A4(new_n346_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n396_), .A2(new_n397_), .B1(new_n324_), .B2(new_n345_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(new_n414_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n413_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n398_), .A2(new_n414_), .A3(new_n346_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n426_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n414_), .A3(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n411_), .A3(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n430_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n431_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n410_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n436_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n434_), .A2(new_n435_), .B1(new_n412_), .B2(new_n411_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT96), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n405_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n401_), .B2(new_n400_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n444_), .A2(new_n406_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n430_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n439_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n395_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT104), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n395_), .A2(KEYINPUT104), .A3(new_n448_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n387_), .A2(new_n205_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n294_), .A2(KEYINPUT27), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n453_), .A2(new_n306_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n392_), .A2(new_n393_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(new_n448_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n452_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(G71gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G99gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n245_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G43gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT85), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT30), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n466_), .B(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n470_), .A2(KEYINPUT86), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(KEYINPUT86), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n309_), .B(KEYINPUT31), .ZN(new_n473_));
  OR3_X1    g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(KEYINPUT86), .A3(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n306_), .A2(new_n453_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n454_), .A2(new_n455_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n448_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT105), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT105), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n456_), .A2(new_n481_), .A3(new_n448_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n476_), .A2(new_n457_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n460_), .A2(new_n476_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT79), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n490_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  OR3_X1    g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n496_), .B(new_n499_), .Z(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n499_), .B(new_n504_), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n496_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n494_), .A2(new_n499_), .A3(new_n495_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n503_), .A2(new_n508_), .A3(new_n512_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n514_), .A2(KEYINPUT81), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT81), .B1(new_n514_), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n485_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT9), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n524_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT64), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(KEYINPUT65), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT64), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n538_), .B(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n543_), .B2(new_n533_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n464_), .A3(new_n536_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n532_), .A2(KEYINPUT67), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(KEYINPUT68), .A3(new_n549_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n529_), .A2(new_n531_), .A3(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n546_), .B1(new_n557_), .B2(new_n523_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G85gat), .B(G92gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT8), .ZN(new_n561_));
  INV_X1    g360(.A(new_n532_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n550_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT66), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT66), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n561_), .B(new_n565_), .C1(new_n562_), .C2(new_n550_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n558_), .A2(new_n559_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n548_), .A2(KEYINPUT68), .A3(new_n549_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT68), .B1(new_n548_), .B2(new_n549_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n529_), .A2(new_n531_), .A3(new_n555_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n555_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n560_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT69), .B1(new_n574_), .B2(new_n546_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n545_), .B1(new_n567_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n579_));
  XOR2_X1   g378(.A(G71gat), .B(G78gat), .Z(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n522_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n564_), .A2(new_n566_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n557_), .A2(new_n523_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n559_), .A3(KEYINPUT8), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n575_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT71), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n567_), .A2(new_n593_), .A3(new_n575_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n545_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n583_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT12), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n584_), .B(new_n587_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G120gat), .B(G148gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT70), .ZN(new_n605_));
  INV_X1    g404(.A(new_n545_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n591_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n596_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n576_), .A2(new_n583_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n605_), .B1(new_n610_), .B2(new_n586_), .ZN(new_n611_));
  AOI211_X1 g410(.A(KEYINPUT70), .B(new_n585_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n598_), .B(new_n604_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n591_), .A2(new_n606_), .A3(new_n583_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n583_), .B1(new_n591_), .B2(new_n606_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n586_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT70), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n610_), .A2(new_n605_), .A3(new_n586_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n604_), .B1(new_n620_), .B2(new_n598_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n521_), .B1(new_n614_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n598_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n603_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n613_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT34), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n576_), .A2(new_n499_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n505_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n595_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n632_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n641_), .B(new_n636_), .C1(new_n595_), .C2(new_n637_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT36), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n642_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n645_), .B(KEYINPUT36), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT76), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT37), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT77), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n594_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n593_), .B1(new_n567_), .B2(new_n575_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n606_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n505_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n641_), .B1(new_n658_), .B2(new_n636_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n642_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n649_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT78), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT37), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT78), .B(new_n649_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n663_), .A2(new_n647_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT77), .B(KEYINPUT37), .C1(new_n648_), .C2(new_n651_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n654_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n496_), .B(new_n583_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G231gat), .A2(G233gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(G127gat), .B(G155gat), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT16), .ZN(new_n673_));
  XNOR2_X1  g472(.A(G183gat), .B(G211gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT17), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT80), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n668_), .A2(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n519_), .A2(new_n631_), .A3(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n487_), .A3(new_n457_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n665_), .A2(new_n647_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n663_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n485_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n681_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n518_), .B1(new_n622_), .B2(new_n626_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G1gat), .B1(new_n694_), .B2(new_n394_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n686_), .A2(new_n695_), .ZN(new_n696_));
  MUX2_X1   g495(.A(new_n686_), .B(new_n696_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g496(.A(new_n456_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n685_), .A2(new_n488_), .A3(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT106), .ZN(new_n700_));
  OAI21_X1  g499(.A(G8gat), .B1(new_n694_), .B2(new_n456_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT39), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n702_), .A3(KEYINPUT40), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1325gat));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  OAI21_X1  g507(.A(G15gat), .B1(new_n694_), .B2(new_n476_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT41), .ZN(new_n710_));
  INV_X1    g509(.A(G15gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n476_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n685_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n685_), .A2(KEYINPUT107), .A3(new_n711_), .A4(new_n712_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n710_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n709_), .A2(KEYINPUT41), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n708_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n715_), .A2(new_n716_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n721_), .A2(KEYINPUT108), .A3(new_n718_), .A4(new_n710_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1326gat));
  OAI21_X1  g522(.A(G22gat), .B1(new_n694_), .B2(new_n448_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT42), .ZN(new_n725_));
  INV_X1    g524(.A(new_n448_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n685_), .A2(new_n415_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1327gat));
  NOR2_X1   g527(.A1(new_n479_), .A2(KEYINPUT105), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n481_), .B1(new_n456_), .B2(new_n448_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n484_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n395_), .A2(KEYINPUT104), .A3(new_n448_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT104), .B1(new_n395_), .B2(new_n448_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n458_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n735_), .B2(new_n712_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n518_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n627_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n688_), .A2(new_n663_), .A3(new_n683_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G29gat), .B1(new_n742_), .B2(new_n457_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n693_), .A2(new_n744_), .A3(new_n683_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n693_), .B2(new_n683_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n654_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n485_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n733_), .A2(new_n734_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n712_), .B1(new_n751_), .B2(new_n452_), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n457_), .B(new_n476_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n750_), .B(new_n668_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n747_), .B1(new_n749_), .B2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(KEYINPUT44), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757_));
  INV_X1    g556(.A(new_n747_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n485_), .A2(KEYINPUT43), .A3(new_n748_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n750_), .B1(new_n736_), .B2(new_n668_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n756_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n457_), .A2(G29gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n743_), .B1(new_n765_), .B2(new_n766_), .ZN(G1328gat));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n456_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n749_), .A2(new_n754_), .ZN(new_n772_));
  AND4_X1   g571(.A1(KEYINPUT110), .A2(new_n772_), .A3(KEYINPUT44), .A4(new_n758_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT110), .B1(new_n755_), .B2(KEYINPUT44), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G36gat), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n456_), .A2(G36gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT45), .B1(new_n741_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n519_), .A2(new_n780_), .A3(new_n740_), .A4(new_n777_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n779_), .A2(new_n781_), .B1(KEYINPUT111), .B2(new_n768_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n770_), .B1(new_n776_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n782_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n769_), .B(new_n784_), .C1(new_n775_), .C2(G36gat), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1329gat));
  AOI21_X1  g585(.A(G43gat), .B1(new_n742_), .B2(new_n712_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n712_), .A2(G43gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n765_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n788_), .B(new_n756_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT47), .B1(new_n793_), .B2(new_n787_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1330gat));
  AOI21_X1  g594(.A(G50gat), .B1(new_n742_), .B2(new_n726_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n448_), .A2(new_n416_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n765_), .B2(new_n797_), .ZN(G1331gat));
  NOR2_X1   g597(.A1(new_n683_), .A2(new_n737_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n691_), .A2(new_n630_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G57gat), .B1(new_n800_), .B2(new_n394_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n485_), .A2(new_n737_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n738_), .A3(new_n684_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n394_), .A2(G57gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(G1332gat));
  OR3_X1    g604(.A1(new_n803_), .A2(G64gat), .A3(new_n456_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n800_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n698_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(G64gat), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(G64gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(G1333gat));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n712_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G71gat), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT49), .B(new_n462_), .C1(new_n807_), .C2(new_n712_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n712_), .A2(new_n462_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n815_), .A2(new_n816_), .B1(new_n803_), .B2(new_n817_), .ZN(G1334gat));
  OR3_X1    g617(.A1(new_n803_), .A2(G78gat), .A3(new_n448_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n807_), .A2(new_n726_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G78gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G78gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(G1335gat));
  NAND3_X1  g623(.A1(new_n738_), .A2(new_n518_), .A3(new_n683_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n749_), .B2(new_n754_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G85gat), .B1(new_n827_), .B2(new_n394_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n739_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(new_n630_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n525_), .A3(new_n457_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1336gat));
  OAI21_X1  g632(.A(G92gat), .B1(new_n827_), .B2(new_n456_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n526_), .A3(new_n698_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n827_), .B2(new_n476_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n712_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n837_), .B(KEYINPUT113), .C1(new_n830_), .C2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g640(.A1(new_n831_), .A2(new_n536_), .A3(new_n726_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n826_), .A2(new_n726_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G106gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT52), .B(new_n536_), .C1(new_n826_), .C2(new_n726_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g647(.A1(new_n483_), .A2(new_n457_), .A3(new_n712_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(new_n683_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n500_), .A2(new_n501_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n506_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n513_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n515_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n614_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n584_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n586_), .B1(new_n858_), .B2(new_n615_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n597_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n657_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT55), .A3(new_n584_), .A4(new_n587_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n598_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(KEYINPUT56), .A3(new_n603_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n865_), .B2(new_n603_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n857_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n748_), .B1(new_n852_), .B2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT58), .B(new_n857_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n518_), .A2(new_n614_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n866_), .B1(new_n868_), .B2(KEYINPUT115), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n874_), .B(KEYINPUT56), .C1(new_n865_), .C2(new_n603_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n872_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n614_), .A2(new_n621_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n856_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n689_), .A2(KEYINPUT57), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n870_), .A2(new_n871_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n865_), .A2(new_n603_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n874_), .B1(new_n885_), .B2(KEYINPUT56), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n868_), .A2(KEYINPUT115), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n866_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n878_), .B1(new_n888_), .B2(new_n872_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n884_), .B1(new_n889_), .B2(new_n690_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n851_), .B1(new_n883_), .B2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n799_), .A2(new_n627_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n892_), .A2(new_n748_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n892_), .B2(new_n748_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n850_), .B1(new_n891_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(G113gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n518_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n869_), .A2(new_n852_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n668_), .A2(new_n900_), .A3(new_n871_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n889_), .B2(new_n881_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n880_), .B2(new_n689_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n681_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n896_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n849_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n897_), .B(new_n899_), .C1(new_n906_), .C2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n905_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n849_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n737_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n898_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n908_), .A2(new_n912_), .A3(KEYINPUT116), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1340gat));
  NOR2_X1   g716(.A1(new_n627_), .A2(KEYINPUT60), .ZN(new_n918_));
  MUX2_X1   g717(.A(new_n918_), .B(KEYINPUT60), .S(G120gat), .Z(new_n919_));
  NAND2_X1  g718(.A1(new_n906_), .A2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT117), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n897_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G120gat), .B1(new_n922_), .B2(new_n631_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1341gat));
  XOR2_X1   g723(.A(KEYINPUT118), .B(G127gat), .Z(new_n925_));
  NOR3_X1   g724(.A1(new_n922_), .A2(new_n681_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G127gat), .B1(new_n906_), .B2(new_n851_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1342gat));
  INV_X1    g727(.A(G134gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n748_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n897_), .B(new_n930_), .C1(new_n906_), .C2(new_n907_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n909_), .A2(new_n690_), .A3(new_n910_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n931_), .A2(new_n933_), .A3(KEYINPUT119), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1343gat));
  AOI21_X1  g737(.A(new_n712_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n698_), .A2(new_n394_), .A3(new_n448_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n518_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n310_), .ZN(G1344gat));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n631_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n311_), .ZN(G1345gat));
  NOR2_X1   g744(.A1(new_n941_), .A2(new_n683_), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT61), .B(G155gat), .Z(new_n947_));
  XNOR2_X1  g746(.A(new_n946_), .B(new_n947_), .ZN(G1346gat));
  OAI21_X1  g747(.A(G162gat), .B1(new_n941_), .B2(new_n748_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n690_), .A2(new_n314_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n941_), .B2(new_n950_), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n891_), .A2(new_n896_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n476_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n726_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(KEYINPUT122), .B1(new_n952_), .B2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n958_), .B(new_n955_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(KEYINPUT22), .B(G169gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n737_), .A2(new_n960_), .ZN(new_n961_));
  XOR2_X1   g760(.A(new_n961_), .B(KEYINPUT123), .Z(new_n962_));
  NAND3_X1  g761(.A1(new_n957_), .A2(new_n959_), .A3(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(G169gat), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n953_), .A2(new_n737_), .ZN(new_n965_));
  OR2_X1    g764(.A1(new_n965_), .A2(KEYINPUT120), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(KEYINPUT120), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n966_), .A2(new_n448_), .A3(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n683_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n905_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT121), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n964_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT121), .B1(new_n952_), .B2(new_n968_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n972_), .A2(new_n973_), .A3(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n974_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n963_), .B1(new_n975_), .B2(new_n976_), .ZN(G1348gat));
  NAND2_X1  g776(.A1(new_n909_), .A2(new_n448_), .ZN(new_n978_));
  INV_X1    g777(.A(G176gat), .ZN(new_n979_));
  NOR4_X1   g778(.A1(new_n978_), .A2(new_n979_), .A3(new_n631_), .A4(new_n954_), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n957_), .A2(new_n738_), .A3(new_n959_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n980_), .B1(new_n979_), .B2(new_n981_), .ZN(G1349gat));
  NOR3_X1   g781(.A1(new_n681_), .A2(new_n235_), .A3(new_n275_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n957_), .A2(new_n959_), .A3(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n953_), .A2(new_n851_), .ZN(new_n985_));
  OAI211_X1 g784(.A(new_n218_), .B(new_n220_), .C1(new_n978_), .C2(new_n985_), .ZN(new_n986_));
  AND2_X1   g785(.A1(new_n984_), .A2(new_n986_), .ZN(G1350gat));
  NAND4_X1  g786(.A1(new_n957_), .A2(new_n690_), .A3(new_n232_), .A4(new_n959_), .ZN(new_n988_));
  AND3_X1   g787(.A1(new_n957_), .A2(new_n668_), .A3(new_n959_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n988_), .B1(new_n989_), .B2(new_n219_), .ZN(G1351gat));
  NAND2_X1  g789(.A1(new_n698_), .A2(new_n458_), .ZN(new_n991_));
  INV_X1    g790(.A(new_n991_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n939_), .A2(new_n992_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n993_), .A2(new_n737_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(KEYINPUT124), .B(G197gat), .ZN(new_n995_));
  INV_X1    g794(.A(new_n995_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n994_), .A2(new_n996_), .ZN(new_n997_));
  NAND3_X1  g796(.A1(new_n993_), .A2(new_n737_), .A3(new_n995_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n997_), .A2(new_n998_), .ZN(G1352gat));
  NAND2_X1  g798(.A1(new_n993_), .A2(new_n630_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n1000_), .A2(G204gat), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n993_), .A2(new_n257_), .A3(new_n630_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1001_), .A2(new_n1002_), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n939_), .A2(new_n692_), .A3(new_n992_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1005_));
  AND2_X1   g804(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1006_));
  NOR3_X1   g805(.A1(new_n1004_), .A2(new_n1005_), .A3(new_n1006_), .ZN(new_n1007_));
  AOI21_X1  g806(.A(new_n1007_), .B1(new_n1004_), .B2(new_n1005_), .ZN(G1354gat));
  NAND3_X1  g807(.A1(new_n939_), .A2(new_n690_), .A3(new_n992_), .ZN(new_n1009_));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n1010_));
  NAND2_X1  g809(.A1(new_n1009_), .A2(new_n1010_), .ZN(new_n1011_));
  NAND4_X1  g810(.A1(new_n939_), .A2(KEYINPUT125), .A3(new_n690_), .A4(new_n992_), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1011_), .A2(new_n1012_), .ZN(new_n1013_));
  XNOR2_X1  g812(.A(KEYINPUT126), .B(G218gat), .ZN(new_n1014_));
  NOR2_X1   g813(.A1(new_n748_), .A2(new_n1014_), .ZN(new_n1015_));
  XOR2_X1   g814(.A(new_n1015_), .B(KEYINPUT127), .Z(new_n1016_));
  AOI22_X1  g815(.A1(new_n1013_), .A2(new_n1014_), .B1(new_n993_), .B2(new_n1016_), .ZN(G1355gat));
endmodule


