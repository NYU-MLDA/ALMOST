//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT68), .B(G71gat), .ZN(new_n206_));
  INV_X1    g005(.A(G78gat), .ZN(new_n207_));
  AOI22_X1  g006(.A1(new_n202_), .A2(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n206_), .A2(new_n207_), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n204_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT69), .ZN(new_n215_));
  INV_X1    g014(.A(new_n204_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n229_));
  OAI22_X1  g028(.A1(new_n228_), .A2(new_n229_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n225_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT6), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G85gat), .B(G92gat), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n237_), .A3(new_n225_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n239_), .A2(KEYINPUT9), .B1(new_n234_), .B2(new_n236_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G106gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT65), .B(G92gat), .ZN(new_n249_));
  INV_X1    g048(.A(G85gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT9), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n247_), .A2(new_n248_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n244_), .A2(new_n245_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n219_), .B(new_n254_), .Z(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n254_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n259_), .A2(new_n260_), .B1(new_n263_), .B2(new_n219_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(KEYINPUT12), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n266_), .A3(new_n256_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G120gat), .B(G148gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(G176gat), .B(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n258_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n258_), .B2(new_n267_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT13), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT78), .B(G8gat), .ZN(new_n283_));
  INV_X1    g082(.A(G1gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G8gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  INV_X1    g089(.A(G36gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G29gat), .ZN(new_n292_));
  INV_X1    g091(.A(G29gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G36gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n292_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n290_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n293_), .A2(G36gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n291_), .A2(G29gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT73), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G43gat), .B(G50gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n289_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n289_), .A2(new_n305_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT81), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n289_), .A2(KEYINPUT81), .A3(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT15), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n296_), .A2(new_n297_), .A3(new_n290_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n303_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n298_), .A2(new_n304_), .A3(KEYINPUT15), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n307_), .B1(new_n318_), .B2(new_n289_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n309_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n322_), .A3(new_n309_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n312_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G113gat), .B(G141gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT83), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT84), .ZN(new_n327_));
  XOR2_X1   g126(.A(G169gat), .B(G197gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n330_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n282_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT95), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT94), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(KEYINPUT94), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(KEYINPUT95), .A3(new_n337_), .A4(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT2), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  OR2_X1    g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n346_), .A2(new_n348_), .B1(new_n349_), .B2(KEYINPUT3), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G155gat), .B(G162gat), .Z(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n345_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(KEYINPUT1), .B2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  XOR2_X1   g161(.A(G127gat), .B(G134gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  AND4_X1   g169(.A1(new_n370_), .A2(new_n353_), .A3(new_n360_), .A4(new_n365_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n359_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n365_), .B1(new_n372_), .B2(new_n370_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND3_X1  g178(.A1(new_n353_), .A2(new_n370_), .A3(new_n360_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n370_), .A3(new_n365_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT99), .B1(new_n384_), .B2(new_n367_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n386_), .B(new_n368_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n375_), .B(new_n379_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n367_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n386_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(KEYINPUT99), .A3(new_n367_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n379_), .B1(new_n393_), .B2(new_n375_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G71gat), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n399_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n400_), .A2(G99gat), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(G99gat), .B1(new_n400_), .B2(new_n401_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G169gat), .A2(G176gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT24), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT89), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT24), .A4(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT23), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G183gat), .A3(G190gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT24), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n417_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n408_), .A2(new_n411_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT86), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT25), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n425_), .B2(G183gat), .ZN(new_n426_));
  INV_X1    g225(.A(G183gat), .ZN(new_n427_));
  AOI211_X1 g226(.A(KEYINPUT87), .B(new_n427_), .C1(new_n422_), .C2(new_n424_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(KEYINPUT85), .A2(G183gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT85), .A2(G183gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(KEYINPUT25), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G190gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT26), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT88), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n432_), .B(new_n435_), .C1(KEYINPUT88), .C2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n419_), .B1(new_n429_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n413_), .A2(new_n415_), .A3(KEYINPUT90), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n412_), .A2(new_n440_), .A3(KEYINPUT23), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(new_n433_), .A3(new_n431_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT91), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n439_), .A2(new_n442_), .A3(new_n445_), .A4(new_n441_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G169gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n438_), .A2(KEYINPUT30), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT30), .B1(new_n438_), .B2(new_n449_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n404_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n411_), .A2(new_n408_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n423_), .A2(KEYINPUT25), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n421_), .A2(KEYINPUT86), .ZN(new_n457_));
  OAI21_X1  g256(.A(G183gat), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT87), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n425_), .A2(new_n420_), .A3(G183gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n437_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n453_), .B1(new_n454_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n398_), .B(G71gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G99gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n438_), .A2(KEYINPUT30), .A3(new_n449_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT92), .B(G43gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT31), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n452_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n452_), .B2(new_n468_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT93), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n470_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n450_), .A2(new_n451_), .A3(new_n404_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n466_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n452_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n473_), .A2(new_n365_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n365_), .B1(new_n473_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n395_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n427_), .A2(new_n433_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n416_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n448_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n409_), .A2(KEYINPUT24), .A3(new_n405_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT25), .B(G183gat), .Z(new_n488_));
  INV_X1    g287(.A(KEYINPUT26), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G190gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n434_), .A2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n487_), .B(new_n418_), .C1(new_n488_), .C2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n439_), .A2(new_n441_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n486_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G197gat), .A2(G204gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(KEYINPUT21), .A3(new_n496_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G211gat), .B(G218gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT20), .B1(new_n494_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT102), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n504_), .B1(new_n454_), .B2(new_n463_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT102), .B(KEYINPUT20), .C1(new_n494_), .C2(new_n504_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G226gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT19), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n504_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n438_), .A2(new_n514_), .A3(new_n449_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n512_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n494_), .B2(new_n504_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G8gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT103), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT103), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT27), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n516_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n514_), .B1(new_n438_), .B2(new_n449_), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT20), .B(new_n516_), .C1(new_n494_), .C2(new_n504_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n534_), .B2(new_n524_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n525_), .A2(new_n528_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n372_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n372_), .B2(new_n539_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G22gat), .B(G50gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n541_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT28), .B1(new_n361_), .B2(KEYINPUT29), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n540_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n537_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n544_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT96), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n504_), .B1(new_n372_), .B2(new_n539_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(G228gat), .A3(G233gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n554_), .B(new_n504_), .C1(new_n372_), .C2(new_n539_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G78gat), .B(G106gat), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n548_), .B(new_n551_), .C1(new_n558_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n545_), .A2(new_n547_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n553_), .A2(KEYINPUT97), .A3(new_n555_), .A4(new_n559_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n530_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n533_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n524_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n524_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n529_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n536_), .A2(new_n568_), .A3(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n483_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n561_), .A2(new_n567_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n536_), .A2(new_n578_), .A3(new_n395_), .A4(new_n575_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n388_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n393_), .A2(KEYINPUT33), .A3(new_n379_), .A4(new_n375_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n571_), .A2(new_n573_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n362_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n366_), .A2(new_n367_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n367_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(new_n379_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n374_), .A2(KEYINPUT101), .A3(new_n367_), .A4(new_n366_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n368_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n379_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT100), .A3(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n587_), .A2(new_n590_), .A3(new_n591_), .A4(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .A4(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n597_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n513_), .A2(new_n519_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(new_n597_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n579_), .B1(new_n602_), .B2(new_n578_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n481_), .A2(new_n482_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n577_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n334_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT34), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT35), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n242_), .A2(new_n253_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(KEYINPUT74), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n244_), .A2(new_n245_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n246_), .A2(new_n252_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n237_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n230_), .A2(new_n225_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(KEYINPUT67), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n240_), .B1(new_n619_), .B2(new_n232_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n317_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT15), .B1(new_n298_), .B2(new_n304_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n616_), .A2(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n609_), .A2(new_n610_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n242_), .A2(new_n253_), .A3(new_n304_), .A4(new_n298_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n623_), .A2(KEYINPUT74), .A3(new_n625_), .A4(new_n611_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT36), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT75), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n628_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n631_), .A2(KEYINPUT36), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n636_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT75), .B(new_n638_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT37), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(KEYINPUT76), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT76), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n627_), .A2(new_n643_), .A3(new_n628_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n632_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n645_), .B(new_n646_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT77), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n641_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n641_), .B2(new_n647_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n289_), .B(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(new_n219_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(new_n261_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n261_), .ZN(new_n656_));
  XOR2_X1   g455(.A(G127gat), .B(G155gat), .Z(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G183gat), .B(G211gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT17), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n655_), .A2(new_n656_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT80), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n661_), .A2(KEYINPUT17), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n654_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n651_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n606_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n395_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n284_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT38), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n637_), .A2(new_n639_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n645_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR4_X1   g479(.A1(new_n334_), .A2(new_n605_), .A3(new_n680_), .A4(new_n669_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n284_), .B1(new_n681_), .B2(new_n673_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n675_), .B2(KEYINPUT38), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n677_), .A2(new_n683_), .ZN(G1324gat));
  OAI21_X1  g483(.A(new_n535_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT103), .B(new_n524_), .C1(new_n513_), .C2(new_n519_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n575_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n672_), .A2(new_n283_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G8gat), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n693_), .B(new_n694_), .Z(G1325gat));
  INV_X1    g494(.A(new_n482_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n473_), .A2(new_n480_), .A3(new_n365_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n397_), .B1(new_n681_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT41), .Z(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT106), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT106), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n672_), .A2(new_n397_), .A3(new_n698_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT107), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n702_), .A3(new_n704_), .ZN(G1326gat));
  INV_X1    g504(.A(G22gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n681_), .B2(new_n578_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT42), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n672_), .A2(new_n706_), .A3(new_n578_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1327gat));
  INV_X1    g509(.A(new_n669_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n679_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n606_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n673_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n669_), .A2(new_n282_), .A3(new_n333_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n395_), .A2(new_n578_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n687_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n578_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n604_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n687_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n698_), .A2(new_n721_), .A3(new_n568_), .A4(new_n395_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n651_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(new_n651_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n716_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  INV_X1    g529(.A(new_n650_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n641_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT43), .B1(new_n605_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n651_), .A3(new_n724_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n715_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n728_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n727_), .A2(KEYINPUT108), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n730_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT44), .B1(new_n727_), .B2(KEYINPUT108), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n737_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT109), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n729_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n395_), .A2(new_n293_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n714_), .B1(new_n744_), .B2(new_n745_), .ZN(G1328gat));
  XOR2_X1   g545(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n747_));
  OAI21_X1  g546(.A(new_n687_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n291_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n721_), .A2(G36gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n713_), .A2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT45), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT45), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n747_), .B1(new_n750_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  INV_X1    g556(.A(new_n748_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n738_), .A2(new_n739_), .A3(new_n730_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT109), .B1(new_n741_), .B2(new_n742_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G36gat), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n757_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n757_), .B(new_n764_), .C1(new_n749_), .C2(new_n291_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n756_), .B1(new_n765_), .B2(new_n767_), .ZN(G1329gat));
  AOI21_X1  g567(.A(G43gat), .B1(new_n713_), .B2(new_n698_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n698_), .A2(G43gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n744_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1330gat));
  INV_X1    g572(.A(G50gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n713_), .A2(new_n774_), .A3(new_n578_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n744_), .A2(new_n776_), .A3(new_n578_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G50gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n744_), .B2(new_n578_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1331gat));
  NOR3_X1   g579(.A1(new_n605_), .A2(new_n333_), .A3(new_n282_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n670_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G57gat), .B1(new_n783_), .B2(new_n673_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT113), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n669_), .A2(new_n282_), .A3(new_n333_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n679_), .A3(new_n723_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT114), .B(G57gat), .Z(new_n788_));
  NOR3_X1   g587(.A1(new_n787_), .A2(new_n395_), .A3(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(new_n789_), .ZN(G1332gat));
  OAI21_X1  g589(.A(G64gat), .B1(new_n787_), .B2(new_n721_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT48), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n721_), .A2(G64gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n782_), .B2(new_n793_), .ZN(G1333gat));
  OAI21_X1  g593(.A(G71gat), .B1(new_n787_), .B2(new_n604_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT49), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n783_), .A2(new_n399_), .A3(new_n698_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1334gat));
  OAI21_X1  g597(.A(G78gat), .B1(new_n787_), .B2(new_n568_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT50), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n783_), .A2(new_n207_), .A3(new_n578_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n734_), .A2(new_n735_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n711_), .A2(new_n333_), .A3(new_n282_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805_), .B2(new_n395_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n781_), .A2(new_n712_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n250_), .A3(new_n673_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1336gat));
  AOI21_X1  g608(.A(G92gat), .B1(new_n807_), .B2(new_n687_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n805_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n687_), .A2(new_n249_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(G1337gat));
  AOI21_X1  g612(.A(new_n222_), .B1(new_n811_), .B2(new_n698_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n698_), .A2(new_n247_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n807_), .B2(new_n815_), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g616(.A1(new_n803_), .A2(new_n578_), .A3(new_n804_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT115), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G106gat), .B1(new_n818_), .B2(KEYINPUT115), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n818_), .A2(KEYINPUT115), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(G106gat), .A4(new_n819_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n807_), .A2(new_n248_), .A3(new_n578_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n256_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n267_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n264_), .A2(new_n266_), .A3(KEYINPUT55), .A4(new_n256_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n272_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT56), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(new_n840_), .A3(new_n272_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n839_), .A2(new_n333_), .A3(new_n274_), .A4(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n324_), .A2(new_n330_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n329_), .B1(new_n319_), .B2(new_n310_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n276_), .B2(new_n275_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n832_), .B1(new_n848_), .B2(new_n680_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n275_), .B1(new_n838_), .B2(KEYINPUT56), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n846_), .A3(new_n841_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n846_), .A4(new_n841_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n651_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n680_), .B1(new_n842_), .B2(new_n847_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT57), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n849_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n669_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n281_), .A2(new_n333_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n711_), .A2(new_n860_), .A3(new_n733_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT54), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n670_), .A2(new_n863_), .A3(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n859_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n576_), .A2(new_n604_), .A3(new_n395_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT59), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n858_), .A2(new_n669_), .B1(new_n864_), .B2(new_n862_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(new_n867_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n831_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n856_), .B(new_n832_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n711_), .B1(new_n874_), .B2(new_n855_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n865_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n333_), .B(new_n867_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(KEYINPUT116), .A3(new_n830_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT116), .B1(new_n877_), .B2(new_n830_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n873_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n873_), .B(KEYINPUT117), .C1(new_n878_), .C2(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1340gat));
  NAND2_X1  g683(.A1(new_n866_), .A2(new_n867_), .ZN(new_n885_));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n282_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(KEYINPUT60), .B2(new_n886_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n885_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n866_), .A2(KEYINPUT59), .A3(new_n867_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n282_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n889_), .B1(new_n892_), .B2(new_n886_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT118), .B(new_n889_), .C1(new_n892_), .C2(new_n886_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1341gat));
  NOR2_X1   g696(.A1(new_n885_), .A2(new_n669_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G127gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n890_), .A2(new_n891_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n711_), .A2(G127gat), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT119), .Z(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(G1342gat));
  INV_X1    g702(.A(G134gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n885_), .B2(new_n679_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT120), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n904_), .B(new_n733_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n604_), .A2(new_n578_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(new_n395_), .A3(new_n687_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n866_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n333_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(G141gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n281_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g716(.A1(new_n911_), .A2(new_n669_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT61), .B(G155gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  OR3_X1    g719(.A1(new_n911_), .A2(G162gat), .A3(new_n679_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G162gat), .B1(new_n911_), .B2(new_n733_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1347gat));
  NAND3_X1  g722(.A1(new_n698_), .A2(new_n395_), .A3(new_n687_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT122), .Z(new_n925_));
  NOR3_X1   g724(.A1(new_n869_), .A2(new_n578_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n333_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n927_), .A2(G169gat), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(G169gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n926_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT22), .B(G169gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n333_), .A2(new_n932_), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(KEYINPUT124), .Z(new_n934_));
  OAI22_X1  g733(.A1(new_n929_), .A2(new_n930_), .B1(new_n931_), .B2(new_n934_), .ZN(G1348gat));
  NAND2_X1  g734(.A1(new_n926_), .A2(new_n281_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G176gat), .ZN(G1349gat));
  OAI211_X1 g736(.A(new_n430_), .B(new_n431_), .C1(new_n931_), .C2(new_n669_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n926_), .A2(new_n711_), .A3(new_n488_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n931_), .B2(new_n733_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n926_), .A2(new_n680_), .A3(new_n436_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n909_), .A2(new_n673_), .A3(new_n721_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n866_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n333_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n281_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n669_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT125), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n945_), .A2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  XOR2_X1   g752(.A(new_n952_), .B(new_n953_), .Z(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n866_), .A2(new_n955_), .A3(new_n680_), .A4(new_n944_), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n866_), .A2(new_n651_), .A3(new_n944_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n955_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(KEYINPUT126), .ZN(G1355gat));
endmodule


