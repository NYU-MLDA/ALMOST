//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(G169gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(G183gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n206_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(G183gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n216_), .B(new_n221_), .C1(new_n226_), .C2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n210_), .A2(KEYINPUT84), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n236_), .A2(new_n209_), .A3(G183gat), .A4(G190gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n208_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n241_), .A2(new_n230_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n216_), .B1(new_n242_), .B2(new_n221_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n215_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(G15gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G71gat), .ZN(new_n249_));
  INV_X1    g048(.A(G99gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n251_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT85), .B(G43gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT31), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n257_), .A2(KEYINPUT86), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n253_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n260_), .B1(new_n263_), .B2(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n205_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT86), .B1(new_n257_), .B2(new_n258_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n260_), .A3(new_n256_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n204_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G218gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G211gat), .ZN(new_n271_));
  INV_X1    g070(.A(G211gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G218gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT91), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT90), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT21), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT21), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT92), .ZN(new_n290_));
  AND2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n281_), .A2(KEYINPUT92), .A3(new_n282_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT21), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n278_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT21), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n271_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n276_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT93), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n289_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n244_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT94), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT19), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n214_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT96), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT96), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n214_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n206_), .A2(KEYINPUT25), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n241_), .A2(new_n230_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n234_), .A2(new_n211_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n234_), .B2(new_n211_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n221_), .B(new_n318_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n303_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n325_), .B(KEYINPUT20), .C1(new_n303_), .C2(new_n244_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n305_), .A2(new_n308_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT101), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n326_), .A2(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT101), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n308_), .A4(new_n305_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n303_), .B2(new_n244_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n312_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n333_), .B1(new_n303_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n307_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT32), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n347_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n348_));
  OR2_X1    g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT87), .B1(new_n347_), .B2(KEYINPUT1), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NOR4_X1   g160(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n353_), .B2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n359_), .B(new_n361_), .C1(new_n362_), .C2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n349_), .A2(new_n347_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n356_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n204_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n205_), .B(new_n356_), .C1(new_n370_), .C2(new_n369_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT4), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n375_), .A3(new_n204_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n346_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n346_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n383_));
  OR3_X1    g182(.A1(new_n377_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n381_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n323_), .A2(new_n303_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(new_n307_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n333_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT97), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n326_), .A2(new_n324_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n243_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n310_), .A2(new_n233_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n232_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n296_), .B1(new_n278_), .B2(new_n295_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT93), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n394_), .A2(new_n397_), .A3(new_n289_), .A4(new_n215_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n325_), .B1(new_n398_), .B2(KEYINPUT20), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n390_), .B(new_n307_), .C1(new_n391_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n305_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n402_), .B2(new_n307_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n389_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n345_), .B(new_n386_), .C1(new_n404_), .C2(new_n344_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n342_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n343_), .B(new_n389_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n385_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT99), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n385_), .A2(new_n409_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT99), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n385_), .A2(new_n413_), .A3(new_n409_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n374_), .A2(new_n346_), .A3(new_n376_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n372_), .A2(new_n373_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n381_), .B1(new_n418_), .B2(new_n382_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .A4(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n408_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n371_), .A2(KEYINPUT29), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT28), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(KEYINPUT28), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n303_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n371_), .B2(KEYINPUT29), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n430_), .A3(new_n425_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(G78gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G22gat), .B(G50gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n429_), .A2(new_n431_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n422_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  INV_X1    g242(.A(new_n389_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n307_), .B1(new_n391_), .B2(new_n399_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT97), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n400_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(new_n343_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n407_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n443_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n441_), .A2(new_n386_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n407_), .A2(KEYINPUT103), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT103), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n447_), .B2(new_n343_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n327_), .A2(KEYINPUT101), .B1(new_n307_), .B2(new_n335_), .ZN(new_n456_));
  AOI211_X1 g255(.A(KEYINPUT102), .B(new_n343_), .C1(new_n456_), .C2(new_n331_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT102), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT27), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n450_), .B(new_n451_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n269_), .B1(new_n442_), .B2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n441_), .B(new_n450_), .C1(new_n455_), .C2(new_n460_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n386_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n269_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT76), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT77), .B(KEYINPUT15), .Z(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  XOR2_X1   g272(.A(G85gat), .B(G92gat), .Z(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT6), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n250_), .A2(new_n435_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(KEYINPUT7), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT67), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n474_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(KEYINPUT68), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n482_), .A2(new_n484_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT66), .B(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  AND2_X1   g287(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n489_));
  OAI22_X1  g288(.A1(KEYINPUT65), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n487_), .A2(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT10), .B(G99gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n476_), .B1(G106gat), .B2(new_n494_), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n485_), .A2(new_n486_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n473_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n493_), .A2(new_n495_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n482_), .A2(new_n484_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n482_), .A2(new_n484_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n471_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n497_), .A2(new_n503_), .A3(new_n504_), .A4(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n471_), .B(new_n472_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n509_), .B(new_n504_), .C1(new_n511_), .C2(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n502_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G190gat), .B(G218gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G134gat), .B(G162gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT36), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(KEYINPUT36), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n510_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n467_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT70), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT11), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT69), .B(G71gat), .Z(new_n529_));
  AOI22_X1  g328(.A1(new_n527_), .A2(new_n528_), .B1(new_n529_), .B2(new_n433_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(new_n433_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT72), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n526_), .A2(new_n532_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n526_), .A2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542_));
  INV_X1    g341(.A(G1gat), .ZN(new_n543_));
  INV_X1    g342(.A(G8gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G1gat), .B(G8gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  AND2_X1   g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  OR2_X1    g349(.A1(new_n541_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT81), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n541_), .A2(new_n550_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n537_), .A2(new_n538_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n550_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n558_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n471_), .A2(new_n548_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n568_), .B(new_n569_), .C1(new_n511_), .C2(new_n548_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n471_), .B(new_n548_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G120gat), .B(G148gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  NAND4_X1  g386(.A1(new_n496_), .A2(new_n535_), .A3(new_n539_), .A4(KEYINPUT12), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n533_), .A2(new_n534_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n508_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT64), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n508_), .A2(new_n589_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(KEYINPUT12), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT12), .B1(new_n496_), .B2(new_n562_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT73), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n591_), .A2(new_n593_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n508_), .A2(KEYINPUT71), .A3(new_n589_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n593_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT71), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n590_), .A2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n600_), .B(new_n601_), .C1(new_n603_), .C2(new_n595_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n587_), .B1(new_n599_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n604_), .A3(new_n587_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(KEYINPUT75), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT75), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(KEYINPUT13), .A3(new_n610_), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n567_), .B(new_n582_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n523_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n464_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n613_), .A2(new_n614_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n582_), .ZN(new_n620_));
  OAI221_X1 g419(.A(KEYINPUT27), .B1(new_n457_), .B2(new_n459_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n464_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n408_), .B2(new_n443_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n621_), .A2(new_n623_), .B1(new_n422_), .B2(new_n441_), .ZN(new_n624_));
  OAI22_X1  g423(.A1(new_n624_), .A2(new_n269_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n521_), .A2(KEYINPUT78), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n519_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n521_), .A2(KEYINPUT78), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n522_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n567_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n626_), .A2(new_n543_), .A3(new_n635_), .A4(new_n386_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n618_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(new_n618_), .ZN(new_n639_));
  OAI221_X1 g438(.A(new_n617_), .B1(new_n618_), .B2(new_n636_), .C1(new_n638_), .C2(new_n639_), .ZN(G1324gat));
  INV_X1    g439(.A(new_n522_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n621_), .A2(new_n450_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n625_), .A2(new_n641_), .A3(new_n615_), .A4(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(G8gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n643_), .B2(G8gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n626_), .A2(new_n635_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n544_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n645_), .A2(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT106), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  OAI221_X1 g450(.A(new_n651_), .B1(new_n647_), .B2(new_n648_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(new_n269_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n647_), .A2(G15gat), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G15gat), .B1(new_n616_), .B2(new_n657_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n616_), .B2(new_n441_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n441_), .A2(G22gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT107), .ZN(new_n668_));
  OAI22_X1  g467(.A1(new_n665_), .A2(new_n666_), .B1(new_n647_), .B2(new_n668_), .ZN(G1327gat));
  NAND2_X1  g468(.A1(new_n522_), .A2(new_n567_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT109), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n620_), .A2(new_n625_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n620_), .A2(new_n625_), .A3(new_n674_), .A4(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n386_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n630_), .A2(new_n680_), .A3(new_n632_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n633_), .A2(KEYINPUT43), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n684_), .A2(KEYINPUT43), .B1(new_n625_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n567_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n619_), .A2(new_n687_), .A3(new_n582_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n679_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n625_), .B2(new_n683_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n685_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n467_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n688_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n690_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n386_), .A2(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n678_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n695_), .A3(new_n642_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n642_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n673_), .A2(new_n675_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT45), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n673_), .A2(new_n705_), .A3(new_n675_), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n700_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n707_), .A3(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  INV_X1    g511(.A(G43gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n657_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n690_), .A2(new_n695_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n690_), .A2(new_n695_), .A3(new_n717_), .A4(new_n714_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n676_), .B2(new_n657_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1330gat));
  OR3_X1    g524(.A1(new_n676_), .A2(G50gat), .A3(new_n441_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n441_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n690_), .A2(new_n695_), .A3(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT113), .ZN(new_n729_));
  OAI21_X1  g528(.A(G50gat), .B1(new_n728_), .B2(KEYINPUT113), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n613_), .A2(new_n614_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n581_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n523_), .A2(new_n687_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n464_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n625_), .A2(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n635_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n464_), .A2(G57gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  OR3_X1    g538(.A1(new_n737_), .A2(G64gat), .A3(new_n701_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G64gat), .B1(new_n734_), .B2(new_n701_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT48), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT48), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1333gat));
  OR3_X1    g543(.A1(new_n737_), .A2(G71gat), .A3(new_n657_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734_), .B2(new_n657_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT49), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT49), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n734_), .B2(new_n441_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n727_), .A2(new_n433_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n751_), .A2(new_n752_), .B1(new_n737_), .B2(new_n753_), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n736_), .A2(new_n671_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n386_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n686_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n733_), .A2(new_n567_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(KEYINPUT114), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n686_), .B2(new_n759_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n464_), .A2(new_n487_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n757_), .B1(new_n764_), .B2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n736_), .A2(new_n642_), .A3(new_n671_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT115), .A3(new_n488_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT115), .B1(new_n767_), .B2(new_n488_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n761_), .A2(G92gat), .A3(new_n642_), .A4(new_n763_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(KEYINPUT116), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1337gat));
  NAND3_X1  g575(.A1(new_n758_), .A2(new_n269_), .A3(new_n760_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G99gat), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n657_), .A2(new_n494_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n756_), .A2(new_n779_), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OR2_X1    g580(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n756_), .A2(new_n435_), .A3(new_n727_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n727_), .B(new_n760_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n784_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n607_), .A2(new_n581_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT119), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n607_), .A2(new_n581_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n599_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n588_), .B(new_n590_), .C1(new_n597_), .C2(KEYINPUT73), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT55), .A3(new_n593_), .A4(new_n598_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n598_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n601_), .B1(new_n803_), .B2(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n587_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n806_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n795_), .B(new_n797_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n568_), .B(new_n572_), .C1(new_n511_), .C2(new_n548_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n577_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n580_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n608_), .A2(new_n610_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n522_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n607_), .A2(new_n813_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n805_), .A2(new_n806_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n634_), .B1(new_n821_), .B2(KEYINPUT58), .ZN(new_n822_));
  INV_X1    g621(.A(new_n816_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI22_X1  g625(.A1(KEYINPUT57), .A2(new_n815_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n795_), .A2(new_n797_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n814_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n641_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n567_), .B1(new_n827_), .B2(new_n833_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n567_), .A2(new_n581_), .A3(KEYINPUT118), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n567_), .B2(new_n581_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n732_), .A2(new_n633_), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n463_), .A2(new_n657_), .A3(new_n464_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n581_), .ZN(new_n845_));
  OR2_X1    g644(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n840_), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n841_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n582_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n843_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n732_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n843_), .B2(new_n687_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n849_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(G127gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n687_), .A2(KEYINPUT121), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(G127gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n857_), .B1(new_n858_), .B2(new_n862_), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n843_), .A2(new_n864_), .A3(new_n522_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n633_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1343gat));
  NAND4_X1  g666(.A1(new_n701_), .A2(new_n657_), .A3(new_n727_), .A4(new_n386_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT122), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n839_), .B2(new_n834_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n581_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n619_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n687_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n870_), .B2(new_n522_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n683_), .A2(G162gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n870_), .B2(new_n879_), .ZN(G1347gat));
  AOI21_X1  g679(.A(new_n701_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n465_), .A2(new_n727_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n581_), .A3(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT62), .B(G169gat), .C1(new_n883_), .C2(KEYINPUT22), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n881_), .A2(new_n581_), .A3(new_n882_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT22), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n217_), .B1(new_n886_), .B2(new_n885_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n884_), .B1(new_n888_), .B2(new_n889_), .ZN(G1348gat));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n882_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n732_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n218_), .ZN(G1349gat));
  NAND2_X1  g692(.A1(new_n230_), .A2(new_n317_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n881_), .A2(new_n687_), .A3(new_n894_), .A4(new_n882_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n896_));
  INV_X1    g695(.A(new_n891_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n897_), .B2(new_n687_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n891_), .B2(new_n633_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n522_), .A2(new_n241_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n891_), .B2(new_n902_), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n269_), .A2(new_n622_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n633_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n821_), .A2(KEYINPUT58), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n831_), .A2(new_n832_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n815_), .A2(KEYINPUT57), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n687_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n838_), .B(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n642_), .B(new_n904_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n840_), .A2(KEYINPUT124), .A3(new_n642_), .A4(new_n904_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916_), .B2(new_n581_), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n279_), .B(new_n582_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1352gat));
  OR2_X1    g718(.A1(new_n280_), .A2(KEYINPUT125), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT126), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n916_), .B2(new_n619_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n732_), .B(new_n923_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1353gat));
  OR2_X1    g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n916_), .B2(new_n687_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT63), .B(G211gat), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n567_), .B(new_n928_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1354gat));
  NAND2_X1  g729(.A1(new_n916_), .A2(new_n522_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n633_), .A2(new_n270_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT127), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n931_), .A2(new_n270_), .B1(new_n916_), .B2(new_n933_), .ZN(G1355gat));
endmodule


