//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT26), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G190gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT78), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n221_), .A2(new_n217_), .A3(G183gat), .A4(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n218_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n219_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(G183gat), .B2(G190gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n216_), .A2(new_n224_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT81), .B1(new_n237_), .B2(KEYINPUT31), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(KEYINPUT31), .B2(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n233_), .B(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n231_), .A2(new_n232_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G15gat), .B(G43gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT79), .Z(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G71gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G99gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n247_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n233_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n250_), .A2(new_n239_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n239_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255_));
  INV_X1    g054(.A(G141gat), .ZN(new_n256_));
  INV_X1    g055(.A(G148gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n258_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n257_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n266_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n259_), .B(new_n268_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G22gat), .B(G50gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT28), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n274_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G197gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT82), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G197gat), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT21), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(G197gat), .B2(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n284_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G218gat), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n291_), .A2(G211gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(G211gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n283_), .A2(new_n295_), .A3(new_n285_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT82), .B(G197gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n282_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT84), .B(new_n298_), .C1(new_n299_), .C2(new_n282_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT21), .B1(new_n292_), .B2(new_n293_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n297_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G228gat), .ZN(new_n308_));
  INV_X1    g107(.A(G233gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n307_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n277_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n283_), .A2(new_n295_), .A3(new_n285_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n295_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n294_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n300_), .B2(new_n284_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n279_), .A2(new_n281_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n289_), .B1(new_n326_), .B2(G204gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n304_), .B1(new_n327_), .B2(KEYINPUT84), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n323_), .A2(new_n325_), .B1(new_n328_), .B2(new_n302_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n312_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n310_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n307_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n315_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n319_), .A2(new_n320_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n320_), .B1(new_n319_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n318_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT86), .B1(new_n316_), .B2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n274_), .B(new_n276_), .Z(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n334_), .B2(KEYINPUT85), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n319_), .A2(new_n334_), .A3(new_n320_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n254_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n229_), .B1(new_n223_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT89), .B(new_n229_), .C1(new_n223_), .C2(new_n347_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT88), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n210_), .A2(KEYINPUT87), .A3(new_n213_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n215_), .B1(new_n225_), .B2(new_n219_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT87), .B1(new_n210_), .B2(new_n213_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n214_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(KEYINPUT88), .A3(new_n354_), .A4(new_n355_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n307_), .B1(new_n352_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n329_), .B2(new_n230_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n350_), .A2(new_n351_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(new_n329_), .A3(new_n358_), .A4(new_n361_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n215_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n224_), .A2(new_n210_), .A3(new_n213_), .A4(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n227_), .A2(new_n229_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n364_), .B(new_n368_), .C1(new_n374_), .C2(new_n307_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n366_), .A2(new_n368_), .B1(new_n370_), .B2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n346_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n329_), .B2(new_n230_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n348_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n307_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n368_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT95), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n368_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n368_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n363_), .A2(new_n391_), .A3(new_n365_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n381_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n383_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n364_), .B1(new_n374_), .B2(new_n307_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n370_), .A2(new_n391_), .A3(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n381_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n375_), .A2(new_n370_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n307_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n369_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n307_), .B2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n400_), .B(new_n382_), .C1(new_n403_), .C2(new_n391_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n346_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n395_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n237_), .A2(new_n273_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n236_), .A2(new_n272_), .A3(new_n267_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n237_), .A2(new_n273_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT91), .A4(new_n411_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G85gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G57gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n418_), .A3(new_n426_), .A4(new_n419_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n345_), .A2(new_n407_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n430_));
  INV_X1    g229(.A(new_n428_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n337_), .A2(new_n343_), .A3(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n407_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT92), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n427_), .A2(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n427_), .A2(KEYINPUT92), .A3(new_n434_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n408_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n424_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT93), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n410_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n410_), .A2(KEYINPUT94), .A3(new_n411_), .A4(new_n414_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(KEYINPUT93), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .A4(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n405_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n400_), .B(new_n451_), .C1(new_n403_), .C2(new_n391_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n428_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n451_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n393_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n344_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n394_), .A2(new_n383_), .B1(new_n405_), .B2(new_n346_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n337_), .A2(new_n431_), .A3(new_n343_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT96), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n433_), .A2(new_n456_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n254_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n429_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G230gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n309_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT10), .B(G99gat), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(G85gat), .B2(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT65), .B(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT64), .B(G85gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT9), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n476_), .B2(KEYINPUT66), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  INV_X1    g277(.A(new_n475_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n479_), .A2(new_n473_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(KEYINPUT9), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n470_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT67), .B(KEYINPUT6), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n466_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT7), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT8), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n494_), .A3(new_n489_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT68), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n482_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n504_));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n482_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n488_), .A2(new_n494_), .A3(new_n489_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n494_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n499_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT69), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n508_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n464_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519_));
  INV_X1    g318(.A(new_n508_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n498_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT12), .B(new_n520_), .C1(new_n521_), .C2(new_n482_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n463_), .B2(new_n309_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n523_), .B1(new_n500_), .B2(new_n508_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n464_), .B1(new_n500_), .B2(new_n508_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT71), .A4(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT5), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G176gat), .B(G204gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n518_), .A2(new_n527_), .A3(new_n530_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n539_), .A2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT77), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G1gat), .B(G8gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(G15gat), .A2(G22gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G15gat), .A2(G22gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G1gat), .A2(G8gat), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n550_), .A2(new_n551_), .B1(KEYINPUT14), .B2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n549_), .A2(new_n553_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G29gat), .B(G36gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT15), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n549_), .B(new_n553_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n562_), .B(new_n559_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n546_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT77), .A4(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(KEYINPUT76), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT76), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n569_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n462_), .A2(new_n545_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n500_), .A2(new_n559_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n560_), .B1(new_n521_), .B2(new_n482_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n590_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n599_), .B(KEYINPUT36), .Z(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT74), .Z(new_n603_));
  OAI21_X1  g402(.A(new_n601_), .B1(new_n596_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT37), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n508_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n562_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n612_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n612_), .A2(new_n618_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n609_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n584_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n428_), .B(KEYINPUT97), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(G1gat), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT38), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n460_), .A2(new_n461_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n429_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n601_), .A2(new_n607_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT98), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635_));
  INV_X1    g434(.A(new_n633_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n462_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n545_), .A2(new_n583_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n622_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n431_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n629_), .A2(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(new_n625_), .ZN(new_n645_));
  INV_X1    g444(.A(G8gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n407_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n641_), .A2(new_n407_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n646_), .C1(new_n641_), .C2(new_n407_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n642_), .B2(new_n461_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n461_), .A2(G15gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n625_), .B2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n344_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n641_), .B2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT42), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n645_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n633_), .A2(new_n622_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n584_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n428_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n605_), .A2(new_n608_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n462_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT101), .B(KEYINPUT43), .C1(new_n670_), .C2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n639_), .A2(new_n623_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n632_), .A2(new_n609_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(KEYINPUT100), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n462_), .B2(new_n669_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n672_), .B(new_n674_), .C1(new_n677_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT43), .B1(new_n676_), .B2(new_n675_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT101), .B1(new_n670_), .B2(new_n671_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n672_), .A4(new_n674_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n626_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n668_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n683_), .A2(new_n407_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n457_), .A2(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n584_), .A2(new_n665_), .A3(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT45), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT102), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n692_), .B2(G36gat), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(KEYINPUT46), .ZN(new_n703_));
  AND4_X1   g502(.A1(KEYINPUT103), .A2(new_n693_), .A3(KEYINPUT46), .A4(new_n697_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT103), .B1(new_n701_), .B2(KEYINPUT46), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n700_), .A2(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(G1329gat));
  INV_X1    g505(.A(G43gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n461_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n689_), .A2(KEYINPUT104), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710_));
  INV_X1    g509(.A(new_n708_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n688_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n666_), .B2(new_n461_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n709_), .A2(new_n716_), .A3(new_n712_), .A4(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  NAND3_X1  g517(.A1(new_n689_), .A2(G50gat), .A3(new_n660_), .ZN(new_n719_));
  INV_X1    g518(.A(G50gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n666_), .B2(new_n344_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT105), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n724_), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n545_), .A2(new_n583_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n623_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT107), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT107), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n431_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT108), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n730_), .A2(new_n736_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n624_), .B2(new_n545_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n582_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n624_), .A2(KEYINPUT106), .A3(new_n545_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n632_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n732_), .B1(new_n741_), .B2(new_n627_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n737_), .A3(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT109), .ZN(G1332gat));
  OR3_X1    g543(.A1(new_n741_), .A2(G64gat), .A3(new_n457_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n730_), .A2(new_n407_), .A3(new_n731_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  OR3_X1    g549(.A1(new_n741_), .A2(G71gat), .A3(new_n461_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n730_), .A2(new_n254_), .A3(new_n731_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(G71gat), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  OR3_X1    g555(.A1(new_n741_), .A2(G78gat), .A3(new_n344_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n730_), .A2(new_n660_), .A3(new_n731_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G78gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G78gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT111), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n727_), .A2(new_n622_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n686_), .A2(new_n672_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n428_), .A2(new_n475_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n727_), .A2(new_n633_), .A3(new_n622_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n632_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n627_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n768_), .A2(new_n769_), .B1(G85gat), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT112), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n768_), .A2(new_n473_), .A3(new_n457_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n771_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G92gat), .B1(new_n776_), .B2(new_n407_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n768_), .B2(new_n461_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n461_), .A2(new_n468_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n771_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(KEYINPUT113), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n781_), .B(new_n783_), .ZN(G1338gat));
  OR3_X1    g583(.A1(new_n771_), .A2(G106gat), .A3(new_n344_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n686_), .A2(new_n660_), .A3(new_n672_), .A4(new_n767_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G106gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G106gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n626_), .A2(new_n457_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n345_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n582_), .A2(new_n538_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n525_), .A2(new_n526_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n528_), .A2(new_n509_), .A3(new_n515_), .A4(new_n522_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n797_), .A2(KEYINPUT55), .B1(new_n798_), .B2(new_n464_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n527_), .A2(new_n800_), .A3(new_n530_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n535_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n796_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n564_), .A2(new_n568_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n573_), .B1(new_n567_), .B2(new_n565_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n575_), .A2(new_n576_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n539_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT57), .B(new_n633_), .C1(new_n807_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT117), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n582_), .A2(new_n538_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n535_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n804_), .B(new_n537_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n636_), .B1(new_n818_), .B2(new_n811_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n810_), .A2(new_n538_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT116), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n805_), .A2(new_n806_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT58), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n609_), .A3(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n822_), .B(new_n830_), .C1(KEYINPUT57), .C2(new_n819_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n623_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n609_), .A2(new_n582_), .A3(new_n623_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  INV_X1    g633(.A(new_n545_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n793_), .B(new_n795_), .C1(new_n832_), .C2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n795_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n633_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(KEYINPUT115), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n822_), .A3(new_n830_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n846_), .A2(new_n822_), .A3(KEYINPUT118), .A4(new_n830_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n623_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n838_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n840_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n839_), .B1(new_n853_), .B2(new_n793_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n583_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n622_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n838_), .B1(new_n858_), .B2(new_n850_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n859_), .B2(new_n840_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n583_), .A2(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n862_), .ZN(G1340gat));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n835_), .B2(KEYINPUT60), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n864_), .A2(KEYINPUT60), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n857_), .A2(new_n860_), .A3(new_n865_), .A4(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n839_), .B(new_n545_), .C1(new_n853_), .C2(new_n793_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(new_n864_), .ZN(G1341gat));
  OAI21_X1  g669(.A(G127gat), .B1(new_n854_), .B2(new_n623_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n623_), .A2(G127gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n857_), .A2(new_n860_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1342gat));
  OAI21_X1  g673(.A(G134gat), .B1(new_n854_), .B2(new_n669_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n633_), .A2(G134gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n857_), .A2(new_n860_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1343gat));
  NOR3_X1   g677(.A1(new_n794_), .A2(new_n254_), .A3(new_n344_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n582_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n545_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n881_), .B2(new_n622_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n859_), .A2(KEYINPUT120), .A3(new_n623_), .A4(new_n880_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n851_), .A2(new_n852_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n622_), .A3(new_n879_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT120), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n881_), .A2(new_n888_), .A3(new_n622_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n886_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n896_), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n881_), .B2(new_n636_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n609_), .A2(G162gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT121), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n881_), .B2(new_n900_), .ZN(G1347gat));
  NAND3_X1  g700(.A1(new_n627_), .A2(new_n254_), .A3(new_n407_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT122), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n344_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT124), .B(new_n905_), .C1(new_n832_), .C2(new_n838_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n838_), .B1(new_n831_), .B2(new_n623_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n904_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT22), .B(G169gat), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n906_), .A2(new_n582_), .A3(new_n909_), .A4(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n903_), .A2(new_n582_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n344_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n913_), .B2(new_n912_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G169gat), .B1(new_n908_), .B2(new_n916_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n911_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n906_), .A2(new_n545_), .A3(new_n909_), .ZN(new_n922_));
  INV_X1    g721(.A(G176gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n835_), .A2(new_n923_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n892_), .A2(new_n905_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n859_), .A2(new_n904_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n929_), .A3(new_n925_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n924_), .A2(new_n927_), .A3(new_n930_), .ZN(G1349gat));
  NAND2_X1  g730(.A1(new_n203_), .A2(new_n205_), .ZN(new_n932_));
  AND4_X1   g731(.A1(new_n932_), .A2(new_n906_), .A3(new_n622_), .A4(new_n909_), .ZN(new_n933_));
  AOI21_X1  g732(.A(G183gat), .B1(new_n928_), .B2(new_n622_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1350gat));
  AND2_X1   g734(.A1(new_n207_), .A2(new_n209_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n906_), .A2(new_n636_), .A3(new_n909_), .A4(new_n936_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n906_), .A2(new_n609_), .A3(new_n909_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n206_), .ZN(G1351gat));
  NOR2_X1   g738(.A1(new_n254_), .A2(new_n344_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n940_), .A2(new_n431_), .A3(new_n407_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n859_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n582_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n545_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g745(.A(new_n941_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n892_), .A2(new_n947_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT63), .B(G211gat), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n948_), .A2(new_n623_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n942_), .A2(new_n622_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  NOR3_X1   g752(.A1(new_n948_), .A2(new_n291_), .A3(new_n669_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n859_), .A2(new_n633_), .A3(new_n941_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956_));
  AOI21_X1  g755(.A(G218gat), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT126), .B1(new_n948_), .B2(new_n633_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n954_), .B1(new_n957_), .B2(new_n958_), .ZN(G1355gat));
endmodule


