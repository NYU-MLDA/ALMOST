//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G141gat), .B(G148gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT94), .ZN(new_n212_));
  NOR3_X1   g011(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT95), .ZN(new_n214_));
  AND2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221_));
  AOI21_X1  g020(.A(new_n212_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G22gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT97), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n224_), .B(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n229_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT98), .B(G197gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G204gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(G197gat), .B2(G204gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(G197gat), .B2(G204gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n235_), .B2(G204gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT99), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n237_), .A2(new_n238_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G228gat), .A3(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT100), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n248_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n254_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n234_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT101), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n250_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n257_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT102), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT102), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(new_n257_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n234_), .A2(new_n255_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n259_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT104), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT103), .B(KEYINPUT18), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT89), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT23), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(KEYINPUT91), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT22), .B(G169gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT90), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT22), .ZN(new_n296_));
  AOI21_X1  g095(.A(G176gat), .B1(new_n296_), .B2(KEYINPUT90), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n290_), .A3(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n291_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(KEYINPUT24), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n279_), .A2(new_n281_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n277_), .A2(KEYINPUT23), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n299_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n248_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n244_), .A2(new_n247_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(new_n286_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n292_), .B1(new_n293_), .B2(new_n303_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n319_), .A2(new_n320_), .B1(new_n283_), .B2(new_n307_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n313_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n299_), .A3(new_n311_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n320_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n283_), .A2(new_n307_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n317_), .B1(new_n327_), .B2(new_n248_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n316_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n276_), .B1(new_n323_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT105), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n315_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n276_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n313_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  OAI211_X1 g137(.A(KEYINPUT105), .B(new_n276_), .C1(new_n323_), .C2(new_n329_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n332_), .A2(new_n315_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n316_), .B1(new_n313_), .B2(new_n322_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT27), .B(new_n336_), .C1(new_n343_), .C2(new_n334_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n270_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347_));
  INV_X1    g146(.A(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT30), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n312_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT92), .B(G15gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT93), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G113gat), .B(G120gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n353_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n211_), .B(KEYINPUT94), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n220_), .A2(new_n221_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n357_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT106), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n366_), .A2(KEYINPUT106), .A3(KEYINPUT4), .A4(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT107), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n366_), .A2(new_n373_), .A3(KEYINPUT4), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(new_n366_), .B2(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n366_), .A2(new_n367_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G57gat), .B(G85gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT109), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G1gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT108), .B(KEYINPUT0), .ZN(new_n386_));
  INV_X1    g185(.A(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n385_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n379_), .A2(new_n381_), .A3(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n361_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n346_), .A2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n269_), .A2(new_n393_), .A3(new_n345_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n372_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n389_), .B1(new_n380_), .B2(new_n378_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n337_), .A2(new_n339_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n379_), .A2(KEYINPUT33), .A3(new_n381_), .A4(new_n389_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT110), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT110), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n399_), .A2(new_n401_), .A3(new_n405_), .A4(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n343_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n323_), .A2(new_n329_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n407_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT111), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(KEYINPUT111), .A3(new_n407_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n393_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n404_), .A2(new_n406_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n396_), .B1(new_n416_), .B2(new_n269_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n361_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n395_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G29gat), .B(G36gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G43gat), .B(G50gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G15gat), .B(G22gat), .ZN(new_n425_));
  INV_X1    g224(.A(G1gat), .ZN(new_n426_));
  INV_X1    g225(.A(G8gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT14), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G8gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n424_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n436_), .B(KEYINPUT88), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n424_), .B(KEYINPUT15), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n431_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n424_), .A2(new_n432_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n434_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G113gat), .B(G141gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G169gat), .B(G197gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  OR2_X1    g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n419_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G232gat), .A2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT34), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT35), .ZN(new_n452_));
  INV_X1    g251(.A(G85gat), .ZN(new_n453_));
  INV_X1    g252(.A(G92gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n455_), .A2(KEYINPUT67), .A3(KEYINPUT9), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n455_), .A2(KEYINPUT67), .A3(new_n456_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT9), .B1(new_n453_), .B2(new_n454_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT64), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT64), .A3(new_n468_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT65), .B(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT66), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n480_), .B(new_n477_), .C1(new_n471_), .C2(new_n475_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n466_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n466_), .B(KEYINPUT68), .C1(new_n479_), .C2(new_n481_), .ZN(new_n485_));
  OR3_X1    g284(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(KEYINPUT69), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n462_), .A2(new_n486_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n455_), .A2(KEYINPUT70), .A3(new_n456_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT8), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT8), .B1(new_n491_), .B2(new_n492_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT73), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n492_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n497_), .B1(new_n500_), .B2(new_n493_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n484_), .B(new_n485_), .C1(new_n496_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n438_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n452_), .B1(new_n503_), .B2(KEYINPUT82), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n494_), .A2(new_n495_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n484_), .A2(new_n424_), .A3(new_n485_), .A4(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n451_), .A2(KEYINPUT35), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT81), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G190gat), .B(G218gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT36), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n508_), .B1(new_n438_), .B2(new_n502_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n438_), .B2(new_n502_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n506_), .B(new_n516_), .C1(new_n518_), .C2(new_n452_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n511_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n514_), .B(KEYINPUT36), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(KEYINPUT84), .A3(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT37), .B1(new_n520_), .B2(new_n523_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT83), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n484_), .A2(new_n485_), .A3(new_n505_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(KEYINPUT11), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT71), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n538_), .A3(KEYINPUT11), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n536_), .B2(KEYINPUT11), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n537_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT71), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n535_), .A4(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT12), .B1(new_n534_), .B2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n542_), .A2(new_n546_), .A3(KEYINPUT74), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT74), .B1(new_n542_), .B2(new_n546_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n502_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n502_), .A2(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT75), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n484_), .A2(new_n505_), .A3(new_n485_), .A4(new_n547_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(KEYINPUT76), .A3(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n556_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n534_), .A2(new_n548_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n559_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n560_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT72), .B(new_n560_), .C1(new_n568_), .C2(new_n559_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n566_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n566_), .B(new_n580_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(KEYINPUT78), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n584_), .A3(new_n578_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n582_), .A2(KEYINPUT79), .A3(new_n583_), .A4(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(KEYINPUT79), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(KEYINPUT79), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT85), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n431_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT86), .Z(new_n594_));
  OR2_X1    g393(.A1(new_n550_), .A2(new_n551_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G127gat), .B(G155gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n595_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT87), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n593_), .B(new_n547_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n600_), .A2(new_n601_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n606_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n533_), .A2(new_n586_), .A3(new_n590_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n449_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n393_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n612_), .A2(G1gat), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n616_));
  INV_X1    g415(.A(new_n524_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n419_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n590_), .A2(new_n586_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n448_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n609_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n426_), .B1(new_n624_), .B2(new_n393_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n615_), .A2(new_n616_), .A3(new_n625_), .ZN(G1324gat));
  XNOR2_X1  g425(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n427_), .B1(new_n624_), .B2(new_n345_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n612_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n427_), .A3(new_n345_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n627_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n628_), .A2(new_n629_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT39), .B(new_n427_), .C1(new_n624_), .C2(new_n345_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n632_), .B(new_n627_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n633_), .A2(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n624_), .B2(new_n418_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(new_n639_), .A3(new_n418_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n624_), .B2(new_n270_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n631_), .A2(new_n644_), .A3(new_n270_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1327gat));
  NAND4_X1  g447(.A1(new_n590_), .A2(new_n448_), .A3(new_n586_), .A4(new_n622_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT113), .Z(new_n650_));
  INV_X1    g449(.A(new_n533_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT114), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n533_), .B2(new_n652_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n419_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n419_), .B2(new_n651_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n650_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n650_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n658_), .A2(G29gat), .A3(new_n393_), .A4(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n609_), .A2(new_n617_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n620_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n449_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n387_), .B1(new_n664_), .B2(new_n613_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n660_), .A2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(new_n345_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n449_), .A2(new_n663_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n449_), .A2(KEYINPUT45), .A3(new_n663_), .A4(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n345_), .A3(new_n659_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G36gat), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(KEYINPUT115), .A3(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(KEYINPUT115), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n676_), .A2(KEYINPUT115), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n675_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1329gat));
  NAND4_X1  g480(.A1(new_n658_), .A2(G43gat), .A3(new_n418_), .A4(new_n659_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n348_), .B1(new_n664_), .B2(new_n361_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1330gat));
  NAND4_X1  g485(.A1(new_n658_), .A2(G50gat), .A3(new_n270_), .A4(new_n659_), .ZN(new_n687_));
  INV_X1    g486(.A(G50gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n664_), .B2(new_n269_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1331gat));
  AND2_X1   g489(.A1(new_n419_), .A2(new_n621_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n622_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n620_), .A3(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT117), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n393_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n619_), .A2(new_n448_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n618_), .A2(new_n609_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n613_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n701_), .A3(new_n345_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n698_), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT48), .B(new_n701_), .C1(new_n703_), .C2(new_n345_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n345_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(G64gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n704_), .B2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n694_), .A2(new_n709_), .A3(new_n418_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT49), .B(new_n709_), .C1(new_n703_), .C2(new_n418_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT49), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n703_), .A2(new_n418_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G71gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n711_), .B2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n694_), .A2(new_n716_), .A3(new_n270_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT50), .B(new_n716_), .C1(new_n703_), .C2(new_n270_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n703_), .A2(new_n270_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n718_), .B2(new_n721_), .ZN(G1335gat));
  AND3_X1   g521(.A1(new_n691_), .A2(new_n620_), .A3(new_n661_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n453_), .A3(new_n393_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n654_), .A2(new_n655_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n619_), .A2(new_n448_), .A3(new_n609_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n393_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n729_), .B2(new_n453_), .ZN(G1336gat));
  NAND3_X1  g529(.A1(new_n723_), .A2(new_n454_), .A3(new_n345_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n345_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(new_n454_), .ZN(G1337gat));
  NAND2_X1  g533(.A1(new_n727_), .A2(new_n418_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G99gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n418_), .A3(new_n476_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT51), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n723_), .A2(new_n270_), .A3(new_n478_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n270_), .B(new_n726_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G106gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G106gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g548(.A(KEYINPUT54), .B1(new_n610_), .B2(new_n448_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n619_), .A2(new_n751_), .A3(new_n621_), .A4(new_n692_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n439_), .A2(new_n440_), .A3(new_n435_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n445_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n442_), .A2(new_n445_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n581_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n549_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n502_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n558_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n559_), .A2(KEYINPUT76), .A3(new_n560_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT76), .B1(new_n559_), .B2(new_n560_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT55), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n556_), .A2(new_n565_), .A3(new_n765_), .A4(new_n558_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n558_), .A2(new_n758_), .A3(new_n759_), .A4(new_n559_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n570_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT118), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n772_), .A3(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n578_), .ZN(new_n775_));
  AOI221_X4 g574(.A(KEYINPUT118), .B1(new_n570_), .B2(new_n768_), .C1(new_n764_), .C2(new_n766_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT56), .B(new_n578_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n757_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n533_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n578_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n778_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT58), .A4(new_n757_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT58), .B(new_n757_), .C1(new_n775_), .C2(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT119), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n782_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n448_), .A2(new_n581_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n785_), .B2(new_n778_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n582_), .A2(new_n756_), .A3(new_n585_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n617_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT57), .B(new_n617_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n753_), .B1(new_n799_), .B2(new_n622_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n346_), .A2(new_n393_), .A3(new_n418_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  OAI22_X1  g603(.A1(new_n800_), .A2(new_n801_), .B1(new_n804_), .B2(KEYINPUT59), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n448_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G113gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n799_), .A2(new_n622_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n753_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n801_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n621_), .A2(G113gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n807_), .B1(new_n812_), .B2(new_n813_), .ZN(G1340gat));
  AND3_X1   g613(.A1(new_n803_), .A2(new_n620_), .A3(new_n805_), .ZN(new_n815_));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n619_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(KEYINPUT60), .B2(new_n816_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n815_), .A2(new_n816_), .B1(new_n812_), .B2(new_n818_), .ZN(G1341gat));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n622_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n805_), .B(new_n821_), .C1(new_n812_), .C2(new_n802_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n812_), .B2(new_n622_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(KEYINPUT121), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT121), .B1(new_n822_), .B2(new_n823_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1342gat));
  NAND3_X1  g625(.A1(new_n803_), .A2(new_n651_), .A3(new_n805_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G134gat), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n617_), .A2(G134gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n812_), .B2(new_n829_), .ZN(G1343gat));
  NOR4_X1   g629(.A1(new_n269_), .A2(new_n418_), .A3(new_n613_), .A4(new_n345_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n810_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n448_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n620_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g636(.A1(new_n832_), .A2(new_n622_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT61), .B(G155gat), .Z(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n832_), .B2(new_n533_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n832_), .A2(G162gat), .A3(new_n617_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n843_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n841_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(G1347gat));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n394_), .A2(new_n269_), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n800_), .A2(new_n667_), .A3(new_n621_), .A4(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G169gat), .B1(new_n851_), .B2(KEYINPUT123), .ZN(new_n852_));
  INV_X1    g651(.A(new_n850_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n810_), .A2(new_n345_), .A3(new_n448_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n851_), .A2(new_n293_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n295_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n851_), .A2(KEYINPUT123), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(KEYINPUT62), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n858_), .A3(new_n861_), .ZN(G1348gat));
  NOR3_X1   g661(.A1(new_n800_), .A2(new_n667_), .A3(new_n850_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n620_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n609_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n300_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n284_), .B2(new_n866_), .ZN(G1350gat));
  NAND2_X1  g667(.A1(new_n524_), .A2(new_n301_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT124), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n863_), .A2(new_n651_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n285_), .ZN(G1351gat));
  NOR2_X1   g672(.A1(new_n800_), .A2(new_n667_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n269_), .A2(new_n418_), .A3(new_n393_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n448_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n620_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g679(.A1(new_n810_), .A2(new_n345_), .A3(new_n609_), .A4(new_n875_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT63), .B(G211gat), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n874_), .A2(new_n609_), .A3(new_n875_), .A4(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1354gat));
  AND3_X1   g687(.A1(new_n874_), .A2(new_n524_), .A3(new_n875_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G218gat), .B1(new_n889_), .B2(KEYINPUT126), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n874_), .A2(new_n875_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n617_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n651_), .A2(G218gat), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n890_), .A2(new_n893_), .B1(new_n876_), .B2(new_n894_), .ZN(G1355gat));
endmodule


