//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_;
  INV_X1    g000(.A(G197gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(new_n202_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n207_), .B2(G204gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n205_), .A2(new_n213_), .A3(new_n206_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n202_), .A2(G204gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n205_), .A2(KEYINPUT85), .A3(new_n213_), .A4(new_n206_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT21), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n212_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT23), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT78), .B(G183gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(G190gat), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n227_), .B(KEYINPUT81), .C1(G190gat), .C2(new_n228_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n234_));
  INV_X1    g033(.A(G169gat), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT22), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT22), .B1(new_n234_), .B2(new_n235_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .A4(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n237_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT24), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n227_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n228_), .B2(KEYINPUT25), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G190gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT26), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n225_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n227_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n237_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n232_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n244_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(KEYINPUT91), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(KEYINPUT91), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n253_), .B1(new_n225_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n252_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n225_), .A2(new_n251_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT20), .ZN(new_n271_));
  INV_X1    g070(.A(new_n257_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n225_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT88), .B(new_n212_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n271_), .B1(new_n276_), .B2(new_n261_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n269_), .B1(new_n277_), .B2(new_n268_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G8gat), .B(G36gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n268_), .B1(new_n252_), .B2(new_n265_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n268_), .B1(new_n225_), .B2(new_n264_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n271_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(KEYINPUT27), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT1), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n292_), .B(KEYINPUT82), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(KEYINPUT83), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT2), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n302_), .B(KEYINPUT3), .Z(new_n307_));
  OAI211_X1 g106(.A(new_n294_), .B(new_n299_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310_));
  INV_X1    g109(.A(G113gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G120gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G120gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n312_), .B(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(new_n308_), .A3(new_n304_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n317_), .A3(KEYINPUT4), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT93), .Z(new_n320_));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n309_), .A2(new_n321_), .A3(new_n313_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G1gat), .B(G29gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(G57gat), .B(G85gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n323_), .A2(new_n325_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n271_), .A2(new_n288_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n284_), .B1(new_n286_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n290_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n291_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n274_), .A2(new_n341_), .A3(new_n275_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n225_), .A2(new_n343_), .A3(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT87), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n225_), .A2(KEYINPUT87), .A3(new_n341_), .A4(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G78gat), .B(G106gat), .Z(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT89), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G22gat), .B(G50gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT28), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n345_), .B(new_n350_), .C1(KEYINPUT89), .C2(new_n352_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT90), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n354_), .A2(new_n362_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n351_), .A2(new_n352_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n351_), .A2(new_n352_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n251_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(new_n313_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT31), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n370_), .B(new_n316_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n368_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(new_n361_), .A3(new_n363_), .A4(new_n367_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n340_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n332_), .A2(KEYINPUT33), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n318_), .A2(new_n324_), .A3(new_n322_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n314_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n330_), .A3(new_n392_), .ZN(new_n393_));
  AND4_X1   g192(.A1(new_n290_), .A2(new_n336_), .A3(new_n390_), .A4(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n332_), .A2(KEYINPUT33), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n283_), .A2(KEYINPUT32), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n334_), .B1(new_n278_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n287_), .A2(new_n289_), .A3(new_n396_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n394_), .A2(new_n395_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n400_), .A2(new_n368_), .A3(new_n387_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n389_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G22gat), .ZN(new_n403_));
  INV_X1    g202(.A(G1gat), .ZN(new_n404_));
  INV_X1    g203(.A(G8gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT14), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G8gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G231gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G57gat), .B(G64gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n413_), .A2(KEYINPUT11), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(KEYINPUT11), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G71gat), .B(G78gat), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n416_), .A3(KEYINPUT11), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n411_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G183gat), .B(G211gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G155gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT75), .B(G127gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n420_), .B1(new_n429_), .B2(KEYINPUT76), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(KEYINPUT76), .B2(new_n429_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n420_), .B(KEYINPUT77), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n427_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G190gat), .B(G218gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G134gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G162gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT36), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT10), .B(G99gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT64), .ZN(new_n442_));
  OR3_X1    g241(.A1(new_n442_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT6), .ZN(new_n445_));
  INV_X1    g244(.A(G85gat), .ZN(new_n446_));
  INV_X1    g245(.A(G92gat), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT9), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G85gat), .B(G92gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n450_), .B2(KEYINPUT9), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT65), .B1(new_n442_), .B2(G106gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n443_), .A2(new_n445_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT7), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n445_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n450_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n445_), .B(KEYINPUT66), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n449_), .B1(new_n459_), .B2(new_n455_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT70), .B(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT15), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n453_), .A2(new_n466_), .A3(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G232gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT34), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(KEYINPUT35), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT35), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n472_), .A2(KEYINPUT35), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n474_), .A3(new_n475_), .A4(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n440_), .B1(new_n477_), .B2(KEYINPUT71), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT36), .A3(new_n439_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480_));
  INV_X1    g279(.A(new_n440_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n473_), .A2(new_n480_), .A3(new_n481_), .A4(new_n476_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(KEYINPUT72), .A2(KEYINPUT37), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n478_), .A2(new_n479_), .A3(new_n482_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT72), .A2(KEYINPUT37), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT73), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n485_), .B(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n402_), .A2(new_n436_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n419_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n462_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n453_), .A2(new_n419_), .A3(new_n461_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT12), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n462_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G230gat), .ZN(new_n497_));
  INV_X1    g296(.A(G233gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n491_), .A2(new_n502_), .A3(new_n492_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n462_), .A2(KEYINPUT67), .A3(new_n490_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G120gat), .B(G148gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  OR3_X1    g310(.A1(new_n506_), .A2(KEYINPUT69), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT69), .B1(new_n506_), .B2(new_n511_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n506_), .A2(new_n511_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n466_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n409_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n467_), .B2(new_n409_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n466_), .B(new_n409_), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(G229gat), .A3(G233gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n235_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n202_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n530_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n519_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n489_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT95), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n334_), .B(KEYINPUT96), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n404_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT38), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n478_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n402_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT97), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n543_), .A2(new_n435_), .A3(new_n534_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n334_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n540_), .B1(new_n404_), .B2(new_n546_), .ZN(G1324gat));
  NAND2_X1  g346(.A1(new_n291_), .A2(new_n339_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G8gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT39), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n536_), .A2(new_n405_), .A3(new_n548_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT98), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(KEYINPUT40), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(G1325gat));
  OR3_X1    g357(.A1(new_n535_), .A2(G15gat), .A3(new_n385_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n544_), .A2(new_n387_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G15gat), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT99), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT99), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n562_), .A2(KEYINPUT41), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT41), .B1(new_n562_), .B2(new_n563_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n559_), .B1(new_n564_), .B2(new_n565_), .ZN(G1326gat));
  INV_X1    g365(.A(G22gat), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n544_), .B2(new_n368_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT42), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n368_), .A2(new_n567_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT100), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n535_), .B2(new_n571_), .ZN(G1327gat));
  INV_X1    g371(.A(G29gat), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT44), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT101), .ZN(new_n575_));
  INV_X1    g374(.A(new_n533_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n436_), .B(new_n576_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n488_), .B1(new_n389_), .B2(new_n401_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT43), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT43), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n488_), .C1(new_n389_), .C2(new_n401_), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n575_), .B(new_n577_), .C1(new_n579_), .C2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT102), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n577_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n575_), .B1(KEYINPUT102), .B2(KEYINPUT44), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n573_), .B1(new_n589_), .B2(new_n538_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT103), .ZN(new_n591_));
  INV_X1    g390(.A(new_n541_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n402_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n577_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n573_), .A3(new_n545_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(G1328gat));
  INV_X1    g397(.A(G36gat), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n593_), .A2(new_n594_), .A3(new_n599_), .A4(new_n548_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT45), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n386_), .A2(new_n388_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n340_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n401_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n580_), .B1(new_n607_), .B2(new_n488_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n581_), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT101), .B(new_n594_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT44), .B1(new_n610_), .B2(KEYINPUT102), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n548_), .B1(new_n611_), .B2(new_n587_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n602_), .B1(new_n612_), .B2(G36gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT104), .B1(new_n613_), .B2(KEYINPUT46), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT46), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n599_), .B1(new_n589_), .B2(new_n548_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n615_), .B(new_n616_), .C1(new_n617_), .C2(new_n602_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n548_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT46), .B(new_n601_), .C1(new_n621_), .C2(new_n599_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n612_), .A2(G36gat), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n625_), .A2(KEYINPUT105), .A3(KEYINPUT46), .A4(new_n601_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n619_), .A2(new_n627_), .A3(KEYINPUT106), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1329gat));
  INV_X1    g431(.A(new_n589_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G43gat), .B1(new_n633_), .B2(new_n385_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n385_), .A2(G43gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n595_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g436(.A(G50gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n596_), .A2(new_n638_), .A3(new_n368_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n589_), .A2(new_n368_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT107), .Z(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n641_), .B2(new_n638_), .ZN(G1331gat));
  NAND2_X1  g441(.A1(new_n519_), .A2(new_n533_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n543_), .A2(new_n435_), .A3(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(G57gat), .A3(new_n545_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT108), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n489_), .A2(new_n644_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G57gat), .B1(new_n649_), .B2(new_n538_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1332gat));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n645_), .B2(new_n548_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT48), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n649_), .A2(new_n652_), .A3(new_n548_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1333gat));
  INV_X1    g455(.A(G71gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n645_), .B2(new_n387_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT49), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n649_), .A2(new_n657_), .A3(new_n387_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1334gat));
  INV_X1    g460(.A(G78gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n645_), .B2(new_n368_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT50), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n649_), .A2(new_n662_), .A3(new_n368_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1335gat));
  NOR2_X1   g465(.A1(new_n643_), .A2(new_n435_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n593_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n446_), .B1(new_n668_), .B2(new_n537_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT109), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n579_), .A2(new_n581_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n667_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n334_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n670_), .B1(new_n675_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g475(.A(new_n668_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G92gat), .B1(new_n677_), .B2(new_n548_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n673_), .A2(new_n674_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n620_), .A2(new_n447_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT111), .Z(G1337gat));
  NOR3_X1   g481(.A1(new_n668_), .A2(new_n385_), .A3(new_n442_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n673_), .A2(new_n674_), .A3(new_n385_), .ZN(new_n685_));
  INV_X1    g484(.A(G99gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT112), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n684_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g491(.A1(new_n672_), .A2(new_n368_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G106gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT52), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n696_), .A3(G106gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n368_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n668_), .A2(G106gat), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT113), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n704_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT53), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1339gat));
  AND2_X1   g507(.A1(new_n501_), .A2(KEYINPUT55), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n501_), .A2(KEYINPUT55), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n709_), .A2(new_n710_), .B1(new_n500_), .B2(new_n496_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT56), .B1(new_n711_), .B2(new_n511_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n576_), .B(new_n514_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n514_), .A2(new_n516_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n525_), .A2(new_n523_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n522_), .B(KEYINPUT115), .Z(new_n718_));
  OAI211_X1 g517(.A(new_n530_), .B(new_n717_), .C1(new_n718_), .C2(new_n523_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(new_n531_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n541_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT57), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n713_), .A2(new_n725_), .B1(new_n513_), .B2(new_n512_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n711_), .A2(new_n511_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(KEYINPUT116), .A3(new_n712_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n726_), .A2(new_n720_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT58), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(KEYINPUT58), .A3(new_n720_), .A4(new_n730_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n488_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n435_), .B1(new_n724_), .B2(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n517_), .A2(new_n518_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n488_), .A2(new_n436_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n533_), .A4(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n736_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n388_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n548_), .A2(new_n537_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n311_), .B1(new_n746_), .B2(new_n533_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n752_));
  NAND4_X1  g551(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .A4(new_n752_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n311_), .B(new_n533_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n749_), .A2(new_n754_), .ZN(G1340gat));
  NOR2_X1   g554(.A1(new_n315_), .A2(KEYINPUT60), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT60), .ZN(new_n757_));
  AOI21_X1  g556(.A(G120gat), .B1(new_n519_), .B2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n746_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT119), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT119), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n737_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n760_), .A2(new_n761_), .B1(new_n315_), .B2(new_n762_), .ZN(G1341gat));
  INV_X1    g562(.A(new_n746_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G127gat), .B1(new_n764_), .B2(new_n435_), .ZN(new_n765_));
  INV_X1    g564(.A(G127gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n767_), .B2(new_n435_), .ZN(G1342gat));
  AOI21_X1  g567(.A(G134gat), .B1(new_n764_), .B2(new_n541_), .ZN(new_n769_));
  INV_X1    g568(.A(G134gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n488_), .ZN(G1343gat));
  INV_X1    g571(.A(new_n386_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n743_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n745_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n533_), .ZN(new_n776_));
  INV_X1    g575(.A(G141gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1344gat));
  NOR2_X1   g577(.A1(new_n775_), .A2(new_n737_), .ZN(new_n779_));
  INV_X1    g578(.A(G148gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1345gat));
  NOR2_X1   g580(.A1(new_n775_), .A2(new_n436_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(G155gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n782_), .B(new_n784_), .ZN(G1346gat));
  INV_X1    g584(.A(new_n775_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G162gat), .B1(new_n786_), .B2(new_n541_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n488_), .A2(G162gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT121), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n786_), .B2(new_n789_), .ZN(G1347gat));
  NOR2_X1   g589(.A1(new_n620_), .A2(new_n538_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n744_), .B(new_n791_), .C1(new_n736_), .C2(new_n742_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n576_), .A2(new_n255_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT122), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n792_), .A2(new_n533_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G169gat), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n796_), .B(G169gat), .C1(new_n792_), .C2(new_n533_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT123), .B(new_n795_), .C1(new_n798_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1348gat));
  NOR2_X1   g604(.A1(new_n792_), .A2(new_n737_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(new_n237_), .ZN(G1349gat));
  NOR2_X1   g606(.A1(new_n792_), .A2(new_n436_), .ZN(new_n808_));
  MUX2_X1   g607(.A(new_n228_), .B(new_n258_), .S(new_n808_), .Z(G1350gat));
  INV_X1    g608(.A(new_n488_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G190gat), .B1(new_n792_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n541_), .A2(new_n259_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n792_), .B2(new_n812_), .ZN(G1351gat));
  NOR2_X1   g612(.A1(new_n620_), .A2(new_n545_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n743_), .A2(new_n773_), .A3(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n533_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT124), .B(G197gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1352gat));
  NAND3_X1  g617(.A1(new_n774_), .A2(new_n519_), .A3(new_n814_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n821_));
  MUX2_X1   g620(.A(new_n819_), .B(new_n820_), .S(new_n821_), .Z(G1353gat));
  XNOR2_X1  g621(.A(KEYINPUT63), .B(G211gat), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n774_), .A2(new_n435_), .A3(new_n814_), .A4(new_n823_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n815_), .A2(new_n436_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT126), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1354gat));
  XNOR2_X1  g627(.A(KEYINPUT127), .B(G218gat), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n815_), .A2(new_n810_), .A3(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n774_), .A2(new_n541_), .A3(new_n814_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1355gat));
endmodule


