//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_;
  XNOR2_X1  g000(.A(G64gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT90), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G8gat), .B(G36gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G226gat), .A2(G233gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT19), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G197gat), .A2(G204gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT84), .B(G197gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(G204gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT84), .ZN(new_n221_));
  INV_X1    g020(.A(G197gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G204gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n218_), .B1(G197gat), .B2(G204gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n217_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n225_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(G204gat), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n214_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT21), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n220_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT85), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G169gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n238_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(G169gat), .B2(G176gat), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  INV_X1    g049(.A(G176gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT77), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT25), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G183gat), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT26), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT26), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G190gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n243_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n246_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n253_), .A2(new_n262_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n236_), .A2(new_n245_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n252_), .A2(new_n249_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n244_), .B1(new_n246_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n262_), .A2(KEYINPUT76), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT25), .B(G183gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G190gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n271_), .B(new_n253_), .C1(new_n272_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n245_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n269_), .B1(new_n278_), .B2(new_n235_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n213_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n245_), .A2(new_n267_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n269_), .B1(new_n235_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n224_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n218_), .B1(new_n283_), .B2(new_n214_), .ZN(new_n284_));
  INV_X1    g083(.A(G218gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G211gat), .ZN(new_n286_));
  INV_X1    g085(.A(G211gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G218gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n284_), .A2(new_n290_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n277_), .A2(new_n291_), .A3(new_n245_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n282_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(new_n212_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n210_), .B1(new_n280_), .B2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n279_), .B(new_n213_), .C1(new_n235_), .C2(new_n281_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n293_), .B2(new_n212_), .ZN(new_n298_));
  AOI211_X1 g097(.A(KEYINPUT87), .B(new_n213_), .C1(new_n282_), .C2(new_n292_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n209_), .B(new_n296_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT27), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n293_), .A2(new_n212_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT87), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n297_), .A3(new_n212_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n306_), .A2(KEYINPUT91), .A3(new_n209_), .A4(new_n296_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT91), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n210_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT83), .Z(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G141gat), .B(G148gat), .Z(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(new_n323_), .C2(new_n321_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  INV_X1    g126(.A(G141gat), .ZN(new_n328_));
  INV_X1    g127(.A(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n235_), .B(new_n317_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n236_), .B1(KEYINPUT29), .B2(new_n338_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n317_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n344_), .B(new_n341_), .C1(new_n342_), .C2(new_n317_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G22gat), .B(G50gat), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n338_), .A2(KEYINPUT29), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n350_), .A2(new_n352_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n349_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT82), .B1(new_n356_), .B2(new_n358_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n346_), .B(new_n347_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n343_), .A2(KEYINPUT86), .A3(new_n344_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n344_), .A2(KEYINPUT86), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n365_), .B(new_n341_), .C1(new_n342_), .C2(new_n317_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n366_), .A3(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT78), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(new_n278_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G71gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n372_), .B(new_n375_), .Z(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT79), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n380_), .B2(new_n379_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n376_), .B(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n315_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n379_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n338_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n326_), .A3(new_n337_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n338_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n388_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n391_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n387_), .A2(KEYINPUT94), .A3(new_n388_), .A4(new_n390_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT93), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n394_), .A2(new_n397_), .A3(new_n404_), .A4(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n385_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT92), .A4(new_n312_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n407_), .A2(KEYINPUT33), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n407_), .A2(KEYINPUT33), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n396_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n387_), .A2(KEYINPUT95), .A3(new_n388_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n391_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n405_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n421_), .B2(new_n405_), .ZN(new_n426_));
  OAI22_X1  g225(.A1(new_n416_), .A2(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n414_), .A2(new_n415_), .A3(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT32), .B(new_n209_), .C1(new_n280_), .C2(new_n294_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n209_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n306_), .A2(new_n296_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n432_), .A3(new_n408_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n368_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n314_), .A2(new_n368_), .A3(new_n409_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n384_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT97), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT97), .B(new_n384_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n411_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  INV_X1    g241(.A(G8gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G8gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n447_), .B(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(G229gat), .A2(G233gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n450_), .B(KEYINPUT15), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n447_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT75), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G113gat), .B(G141gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G169gat), .B(G197gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n460_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G85gat), .B(G92gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT8), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G57gat), .B(G64gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT11), .ZN(new_n477_));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(KEYINPUT11), .B2(new_n476_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n477_), .A2(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT9), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n466_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(KEYINPUT9), .B2(new_n466_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n485_), .B(KEYINPUT65), .C1(KEYINPUT9), .C2(new_n466_), .ZN(new_n489_));
  INV_X1    g288(.A(G106gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n473_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n475_), .A2(new_n482_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n475_), .A2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n482_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G230gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT64), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(KEYINPUT67), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n475_), .A2(new_n505_), .A3(new_n493_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n504_), .A2(KEYINPUT12), .A3(new_n498_), .A4(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT68), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(new_n507_), .A3(new_n510_), .A4(new_n503_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n499_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n502_), .B1(new_n512_), .B2(new_n495_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G120gat), .B(G148gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT5), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G176gat), .B(G204gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n509_), .A2(new_n511_), .A3(new_n513_), .A4(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(KEYINPUT13), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT13), .B1(new_n519_), .B2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n440_), .A2(new_n465_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n475_), .A2(new_n493_), .A3(new_n450_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n504_), .A2(new_n506_), .A3(new_n455_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n529_), .A2(new_n530_), .A3(new_n539_), .A4(new_n535_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(KEYINPUT71), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n538_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(new_n548_), .A3(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT37), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(KEYINPUT37), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(KEYINPUT37), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n551_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n447_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n498_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT73), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT16), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n562_), .B(new_n567_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n561_), .A2(KEYINPUT17), .A3(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT74), .Z(new_n571_));
  NOR2_X1   g370(.A1(new_n558_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n526_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n442_), .A3(new_n408_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n524_), .A2(KEYINPUT98), .A3(new_n464_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT98), .B1(new_n524_), .B2(new_n464_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n570_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n552_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n439_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n314_), .A2(new_n368_), .A3(new_n409_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n433_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n427_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n586_), .B2(new_n415_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n587_), .B2(new_n368_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT97), .B1(new_n588_), .B2(new_n384_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n410_), .B1(new_n583_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n582_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n409_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n576_), .A2(new_n577_), .A3(new_n592_), .ZN(G1324gat));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n314_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n594_), .A2(KEYINPUT100), .A3(new_n443_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT100), .B1(new_n594_), .B2(new_n443_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT39), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n573_), .A2(new_n443_), .A3(new_n315_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT99), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT100), .B(new_n600_), .C1(new_n594_), .C2(new_n443_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(G1325gat));
  INV_X1    g403(.A(G15gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n384_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n573_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n582_), .A2(new_n606_), .A3(new_n590_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n608_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT41), .B1(new_n608_), .B2(G15gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT102), .Z(G1326gat));
  INV_X1    g411(.A(new_n368_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G22gat), .B1(new_n591_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n573_), .A2(new_n616_), .A3(new_n368_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1327gat));
  INV_X1    g417(.A(new_n571_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n552_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n526_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n622_), .B2(new_n408_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n580_), .B2(new_n619_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT103), .B(new_n571_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n590_), .A2(new_n628_), .A3(new_n629_), .A4(new_n558_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n558_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT43), .B1(new_n440_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n438_), .A2(new_n439_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n631_), .B1(new_n634_), .B2(new_n410_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n628_), .B1(new_n635_), .B2(new_n629_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n627_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT44), .B(new_n627_), .C1(new_n633_), .C2(new_n636_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n408_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n623_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n639_), .A2(new_n315_), .A3(new_n640_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n314_), .A2(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n526_), .A2(new_n621_), .A3(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT45), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n644_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n645_), .B2(G36gat), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n656_));
  AND4_X1   g455(.A1(new_n656_), .A2(new_n646_), .A3(KEYINPUT46), .A4(new_n650_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n654_), .B2(KEYINPUT46), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n653_), .A2(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1329gat));
  NAND3_X1  g458(.A1(new_n641_), .A2(G43gat), .A3(new_n606_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G43gat), .B1(new_n622_), .B2(new_n606_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT107), .Z(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1330gat));
  AOI21_X1  g465(.A(G50gat), .B1(new_n622_), .B2(new_n368_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n368_), .A2(G50gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n641_), .B2(new_n668_), .ZN(G1331gat));
  NOR3_X1   g468(.A1(new_n440_), .A2(new_n464_), .A3(new_n524_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(G57gat), .A3(new_n408_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT110), .Z(new_n673_));
  INV_X1    g472(.A(G57gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n572_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n408_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n673_), .B1(new_n674_), .B2(new_n679_), .ZN(G1332gat));
  NAND2_X1  g479(.A1(new_n671_), .A2(new_n315_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G64gat), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT48), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n314_), .A2(G64gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n675_), .B2(new_n684_), .ZN(G1333gat));
  AOI21_X1  g484(.A(new_n374_), .B1(new_n671_), .B2(new_n606_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT49), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n676_), .A2(new_n374_), .A3(new_n606_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n671_), .B2(new_n368_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT50), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n676_), .A2(new_n690_), .A3(new_n368_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1335gat));
  AND2_X1   g493(.A1(new_n670_), .A2(new_n621_), .ZN(new_n695_));
  INV_X1    g494(.A(G85gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n408_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n633_), .A2(new_n636_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n524_), .A2(new_n464_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n571_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n408_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n697_), .B1(new_n703_), .B2(new_n696_), .ZN(G1336gat));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G92gat), .B1(new_n705_), .B2(new_n314_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n695_), .A2(new_n483_), .A3(new_n315_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1337gat));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n491_), .A3(new_n606_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT111), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n712_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G99gat), .B1(new_n705_), .B2(new_n384_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1338gat));
  NAND3_X1  g518(.A1(new_n695_), .A2(new_n490_), .A3(new_n368_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n701_), .A2(new_n368_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G106gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT52), .B(new_n490_), .C1(new_n701_), .C2(new_n368_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT53), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1339gat));
  NOR2_X1   g528(.A1(new_n525_), .A2(new_n464_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT54), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n572_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n572_), .B2(new_n730_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n509_), .A2(new_n511_), .A3(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT114), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n508_), .A2(new_n737_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n503_), .B1(new_n500_), .B2(new_n507_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n738_), .B2(KEYINPUT114), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n518_), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n521_), .A2(new_n464_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n521_), .A2(KEYINPUT113), .A3(new_n464_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n744_), .A2(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n518_), .B(new_n745_), .C1(new_n739_), .C2(new_n743_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n519_), .A2(new_n521_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n452_), .A2(new_n453_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n463_), .B(new_n754_), .C1(new_n453_), .C2(new_n457_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT116), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n751_), .A2(new_n752_), .B1(new_n753_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n736_), .B1(new_n758_), .B2(new_n552_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n752_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n753_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n552_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT57), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n744_), .A2(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n744_), .A2(KEYINPUT56), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n757_), .A2(new_n521_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(KEYINPUT58), .A3(new_n767_), .A4(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n558_), .A3(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT118), .B(new_n736_), .C1(new_n758_), .C2(new_n552_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n761_), .A2(new_n765_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n734_), .B1(new_n775_), .B2(new_n581_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n385_), .A2(new_n408_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779_), .B2(new_n464_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT59), .B1(new_n776_), .B2(new_n778_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n776_), .C2(new_n778_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n773_), .A2(new_n765_), .A3(new_n759_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n734_), .B1(new_n785_), .B2(new_n571_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n778_), .A2(KEYINPUT59), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT120), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n571_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n734_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n787_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n783_), .A2(new_n784_), .B1(new_n789_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n464_), .A2(G113gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT121), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n780_), .B1(new_n795_), .B2(new_n797_), .ZN(G1340gat));
  INV_X1    g597(.A(G120gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n524_), .B2(KEYINPUT60), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n779_), .B(new_n800_), .C1(KEYINPUT60), .C2(new_n799_), .ZN(new_n801_));
  AOI221_X4 g600(.A(new_n524_), .B1(new_n789_), .B2(new_n794_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n799_), .ZN(G1341gat));
  INV_X1    g602(.A(G127gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n779_), .A2(new_n804_), .A3(new_n619_), .ZN(new_n805_));
  AOI221_X4 g604(.A(new_n581_), .B1(new_n789_), .B2(new_n794_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(G1342gat));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n779_), .A2(new_n808_), .A3(new_n552_), .ZN(new_n809_));
  AOI221_X4 g608(.A(new_n631_), .B1(new_n789_), .B2(new_n794_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1343gat));
  NAND2_X1  g610(.A1(new_n775_), .A2(new_n581_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n791_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n606_), .A2(new_n613_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n408_), .A3(new_n314_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT122), .Z(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(KEYINPUT123), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(KEYINPUT123), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n464_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G141gat), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n328_), .B(new_n464_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1344gat));
  OAI21_X1  g622(.A(new_n525_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G148gat), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n329_), .B(new_n525_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1345gat));
  OAI21_X1  g626(.A(new_n619_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n829_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n619_), .B(new_n831_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1346gat));
  INV_X1    g632(.A(new_n819_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n817_), .A2(KEYINPUT123), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n631_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G162gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n818_), .A2(new_n819_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n552_), .A2(new_n837_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n836_), .A2(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(G1347gat));
  NOR2_X1   g639(.A1(new_n314_), .A2(new_n408_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n606_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n368_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n786_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT22), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n464_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT62), .A3(new_n250_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n786_), .A2(new_n465_), .A3(new_n844_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n846_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n792_), .A2(new_n849_), .A3(new_n464_), .A4(new_n843_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G169gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n848_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT124), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n848_), .B(new_n856_), .C1(new_n851_), .C2(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1348gat));
  AOI21_X1  g657(.A(G176gat), .B1(new_n845_), .B2(new_n525_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n776_), .A2(new_n368_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n524_), .A2(new_n251_), .A3(new_n842_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1349gat));
  NOR2_X1   g661(.A1(new_n571_), .A2(new_n842_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G183gat), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n792_), .A2(new_n843_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n581_), .A3(new_n274_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1350gat));
  OAI21_X1  g668(.A(G190gat), .B1(new_n865_), .B2(new_n631_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n845_), .A2(new_n552_), .A3(new_n275_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1351gat));
  AND2_X1   g671(.A1(new_n814_), .A2(new_n841_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n813_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n465_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n222_), .ZN(G1352gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n524_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n224_), .ZN(G1353gat));
  INV_X1    g677(.A(new_n874_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n570_), .B1(new_n880_), .B2(new_n287_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT126), .Z(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n287_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1354gat));
  INV_X1    g684(.A(KEYINPUT127), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n874_), .A2(new_n631_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n285_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n874_), .A2(G218gat), .A3(new_n620_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n886_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n879_), .A2(new_n285_), .A3(new_n552_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(KEYINPUT127), .C1(new_n285_), .C2(new_n887_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1355gat));
endmodule


