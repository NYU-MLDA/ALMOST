//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G85gat), .B(G92gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT65), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n204_), .B1(new_n207_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT8), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n203_), .B1(KEYINPUT9), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  AOI21_X1  g022(.A(new_n207_), .B1(new_n210_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT34), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT35), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n234_), .A2(KEYINPUT71), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n230_), .B(KEYINPUT15), .Z(new_n236_));
  OAI211_X1 g035(.A(new_n231_), .B(new_n235_), .C1(new_n236_), .C2(new_n227_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(KEYINPUT35), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT70), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G190gat), .B(G218gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G134gat), .B(G162gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT36), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(KEYINPUT36), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n240_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n240_), .A2(new_n244_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT72), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n202_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n202_), .ZN(new_n251_));
  NOR4_X1   g050(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT72), .A4(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT74), .B(G15gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G22gat), .ZN(new_n255_));
  INV_X1    g054(.A(G1gat), .ZN(new_n256_));
  INV_X1    g055(.A(G8gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT14), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G1gat), .B(G8gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G231gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT66), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G71gat), .B(G78gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n264_), .A2(KEYINPUT66), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(KEYINPUT66), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n266_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(KEYINPUT11), .A3(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n263_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G127gat), .B(G155gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT16), .ZN(new_n278_));
  XOR2_X1   g077(.A(G183gat), .B(G211gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n276_), .A2(KEYINPUT17), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(KEYINPUT17), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n282_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n253_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G43gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT30), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT78), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(G169gat), .B2(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT24), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  INV_X1    g103(.A(G183gat), .ZN(new_n305_));
  INV_X1    g104(.A(G190gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(KEYINPUT25), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT77), .B1(new_n305_), .B2(KEYINPUT25), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(G183gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .A4(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT24), .B1(new_n296_), .B2(new_n298_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n303_), .A2(new_n309_), .A3(new_n316_), .A4(new_n318_), .ZN(new_n319_));
  OR3_X1    g118(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n307_), .B(new_n308_), .C1(G183gat), .C2(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n293_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n293_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  INV_X1    g129(.A(G15gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n332_), .A3(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(KEYINPUT79), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT31), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT31), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(KEYINPUT79), .A3(new_n338_), .A4(new_n335_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G134gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT80), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G155gat), .A3(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n355_), .B2(KEYINPUT1), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT81), .B1(new_n362_), .B2(new_n357_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n348_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n346_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n366_), .A2(new_n368_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n357_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n355_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n342_), .B1(new_n364_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n353_), .B1(G155gat), .B2(G162gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n351_), .A2(KEYINPUT80), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT1), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n359_), .A3(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n356_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n363_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n349_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n342_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n373_), .A3(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n375_), .A2(new_n384_), .A3(KEYINPUT90), .A4(KEYINPUT4), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT91), .Z(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n375_), .B2(KEYINPUT4), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n374_), .B1(new_n381_), .B2(new_n349_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(new_n383_), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n342_), .B(new_n374_), .C1(new_n381_), .C2(new_n349_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n391_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT93), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n256_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n403_));
  INV_X1    g202(.A(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n402_), .B(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n394_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n392_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n398_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n345_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(KEYINPUT82), .Z(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT29), .B1(new_n364_), .B2(new_n374_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G197gat), .A2(G204gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(G197gat), .A2(G204gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(KEYINPUT21), .A3(new_n420_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G211gat), .B(G218gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n425_), .A2(new_n426_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(KEYINPUT83), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n417_), .B1(new_n418_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n432_), .B(new_n417_), .C1(new_n395_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n415_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n432_), .B1(new_n395_), .B2(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n417_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n435_), .A3(new_n414_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n395_), .B2(new_n434_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n395_), .A2(new_n442_), .A3(new_n434_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G22gat), .B(G50gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n443_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n437_), .A2(new_n441_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n435_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT85), .B1(new_n452_), .B2(new_n415_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n454_), .B(new_n414_), .C1(new_n440_), .C2(new_n435_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n447_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT84), .B1(new_n433_), .B2(new_n436_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n440_), .A2(new_n459_), .A3(new_n435_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n414_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n451_), .B1(new_n457_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n299_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n314_), .A2(G183gat), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n311_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n310_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n296_), .A3(new_n298_), .A4(new_n301_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n470_), .A2(new_n473_), .A3(new_n474_), .A4(new_n309_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n322_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n320_), .A2(KEYINPUT87), .A3(new_n321_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n324_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n427_), .A2(new_n428_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n427_), .B(new_n428_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n467_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n432_), .A2(new_n326_), .A3(KEYINPUT88), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT88), .B1(new_n432_), .B2(new_n326_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n466_), .B(new_n485_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G64gat), .B(G92gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n432_), .A2(new_n480_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n316_), .A2(new_n309_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n317_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(new_n324_), .B2(new_n323_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n484_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n498_), .A3(KEYINPUT20), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n465_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n488_), .A2(new_n493_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n488_), .B2(new_n500_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n463_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n500_), .A3(new_n493_), .ZN(new_n504_));
  AND4_X1   g303(.A1(KEYINPUT20), .A2(new_n494_), .A3(new_n498_), .A4(new_n466_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n465_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n493_), .B(KEYINPUT97), .Z(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT27), .B(new_n504_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n462_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n413_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n407_), .A2(new_n503_), .A3(new_n509_), .A4(new_n410_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT98), .B1(new_n462_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n437_), .A2(new_n454_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n450_), .A2(new_n447_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n452_), .A2(KEYINPUT85), .A3(new_n415_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n461_), .A2(new_n515_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n451_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n412_), .A2(new_n520_), .A3(new_n510_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n488_), .A2(new_n500_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n493_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n375_), .A2(KEYINPUT95), .A3(new_n384_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n391_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n408_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n391_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n375_), .B2(KEYINPUT4), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n525_), .B(new_n504_), .C1(new_n530_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n409_), .A2(new_n398_), .A3(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n407_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n493_), .A2(KEYINPUT32), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n523_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n506_), .A2(new_n465_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(new_n541_), .C1(new_n544_), .C2(new_n505_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT96), .B1(new_n507_), .B2(new_n540_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n537_), .A2(new_n539_), .B1(new_n547_), .B2(new_n411_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n514_), .B(new_n522_), .C1(new_n548_), .C2(new_n520_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n345_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n512_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n261_), .B(new_n230_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n261_), .A2(new_n236_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n261_), .B2(new_n230_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n552_), .A2(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G113gat), .B(G141gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT76), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n557_), .A2(new_n562_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n551_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(new_n270_), .B(new_n268_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n267_), .B1(new_n265_), .B2(KEYINPUT11), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n272_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n226_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n275_), .A2(new_n215_), .A3(new_n225_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(KEYINPUT12), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n226_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n569_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n568_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT68), .Z(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT69), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(KEYINPUT13), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n290_), .A2(new_n567_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n256_), .A3(new_n411_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT99), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT38), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n551_), .A2(new_n248_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n566_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n593_), .A4(new_n288_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n412_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  INV_X1    g403(.A(new_n510_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n594_), .A2(new_n257_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT100), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n601_), .A2(new_n510_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n257_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT101), .B1(new_n601_), .B2(new_n510_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT39), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT39), .B1(new_n610_), .B2(new_n611_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n604_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(KEYINPUT40), .A3(new_n612_), .A4(new_n607_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n601_), .B2(new_n550_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT41), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n594_), .A2(new_n331_), .A3(new_n345_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n601_), .B2(new_n462_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n594_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n462_), .A2(G22gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT103), .Z(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n626_), .B2(new_n628_), .ZN(G1327gat));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n289_), .A2(new_n630_), .A3(new_n248_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n246_), .A2(new_n247_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT104), .B1(new_n632_), .B2(new_n288_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n590_), .A2(new_n592_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n567_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n411_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n566_), .B(new_n288_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n549_), .A2(new_n550_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n512_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n642_), .B2(new_n253_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n250_), .A2(new_n252_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n551_), .A2(new_n644_), .A3(KEYINPUT43), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n638_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT44), .B(new_n638_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n412_), .A2(new_n404_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n637_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  NOR2_X1   g451(.A1(new_n510_), .A2(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n567_), .A2(new_n634_), .A3(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(KEYINPUT45), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT45), .B1(new_n655_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(new_n605_), .A3(new_n649_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G36gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n659_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND3_X1  g467(.A1(new_n650_), .A2(G43gat), .A3(new_n345_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G43gat), .B1(new_n636_), .B2(new_n345_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n636_), .B2(new_n520_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n520_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n650_), .B2(new_n675_), .ZN(G1331gat));
  AND2_X1   g475(.A1(new_n590_), .A2(new_n592_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n599_), .A2(new_n677_), .A3(new_n566_), .A4(new_n288_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT109), .B(G57gat), .Z(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n412_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n551_), .A2(new_n600_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n290_), .A2(new_n681_), .A3(new_n677_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT107), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n411_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n680_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  OR3_X1    g487(.A1(new_n683_), .A2(G64gat), .A3(new_n510_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G64gat), .B1(new_n678_), .B2(new_n510_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT48), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT48), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT110), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n689_), .B(new_n695_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1333gat));
  OAI21_X1  g496(.A(G71gat), .B1(new_n678_), .B2(new_n550_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT49), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n550_), .A2(G71gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n683_), .B2(new_n700_), .ZN(G1334gat));
  OAI21_X1  g500(.A(G78gat), .B1(new_n678_), .B2(new_n462_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n462_), .A2(G78gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n683_), .B2(new_n704_), .ZN(G1335gat));
  OR2_X1    g504(.A1(new_n643_), .A2(new_n645_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n593_), .A2(new_n600_), .A3(new_n288_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT111), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n412_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n593_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n681_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G85gat), .A3(new_n412_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1336gat));
  OAI21_X1  g513(.A(G92gat), .B1(new_n709_), .B2(new_n510_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n712_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n217_), .A3(new_n605_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1337gat));
  OAI21_X1  g517(.A(G99gat), .B1(new_n708_), .B2(new_n550_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n345_), .A3(new_n223_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(KEYINPUT112), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n721_), .B(new_n723_), .ZN(G1338gat));
  NOR3_X1   g523(.A1(new_n712_), .A2(G106gat), .A3(new_n462_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n520_), .A3(new_n707_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G106gat), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n726_), .A2(new_n734_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  NOR3_X1   g535(.A1(new_n550_), .A2(new_n511_), .A3(new_n412_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n575_), .A2(new_n577_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(KEYINPUT55), .A3(new_n568_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n578_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT114), .B1(new_n739_), .B2(new_n568_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n575_), .A2(new_n746_), .A3(new_n569_), .A4(new_n577_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n739_), .A2(new_n568_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n745_), .A2(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n744_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n744_), .B2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n584_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n584_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n755_), .A2(new_n600_), .A3(new_n586_), .A4(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n552_), .A2(new_n553_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n553_), .B1(new_n261_), .B2(new_n230_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n555_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n561_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n563_), .A2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT117), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n588_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n758_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n738_), .B1(new_n766_), .B2(new_n632_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n248_), .C1(new_n758_), .C2(new_n765_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n755_), .A2(new_n586_), .A3(new_n764_), .A4(new_n757_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n644_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n585_), .B(KEYINPUT68), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n754_), .B2(KEYINPUT56), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n775_), .A2(KEYINPUT58), .A3(new_n764_), .A4(new_n757_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n288_), .B1(new_n770_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n290_), .A2(new_n566_), .A3(new_n593_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n737_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n771_), .A2(new_n772_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n253_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n776_), .A2(KEYINPUT119), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n766_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n248_), .B1(new_n758_), .B2(new_n765_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n738_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n289_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n781_), .B(KEYINPUT54), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT59), .A3(new_n737_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n786_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n600_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n801_), .B2(new_n800_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(new_n600_), .A3(new_n737_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n799_), .A2(new_n803_), .B1(new_n804_), .B2(new_n800_), .ZN(G1340gat));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(KEYINPUT60), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n797_), .A2(new_n737_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n593_), .B1(new_n786_), .B2(new_n798_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n806_), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n797_), .A2(new_n812_), .A3(new_n288_), .A4(new_n737_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n289_), .B1(new_n786_), .B2(new_n798_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1342gat));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(G134gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n644_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n797_), .A2(new_n248_), .A3(new_n737_), .ZN(new_n818_));
  INV_X1    g617(.A(G134gat), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n799_), .A2(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(G1343gat));
  NOR2_X1   g619(.A1(new_n345_), .A2(new_n462_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(new_n605_), .A3(new_n412_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n797_), .A2(new_n600_), .A3(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT122), .B(G141gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1344gat));
  NAND3_X1  g625(.A1(new_n797_), .A2(new_n677_), .A3(new_n823_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n797_), .A2(new_n288_), .A3(new_n823_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  NAND2_X1  g630(.A1(new_n797_), .A2(new_n823_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G162gat), .B1(new_n832_), .B2(new_n644_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n632_), .A2(G162gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(new_n834_), .ZN(G1347gat));
  NAND2_X1  g634(.A1(new_n605_), .A2(new_n462_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n413_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT22), .B(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n600_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT124), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n838_), .B(new_n841_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n838_), .A2(new_n566_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(G169gat), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n842_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n844_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT123), .B1(new_n850_), .B2(new_n294_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n843_), .A3(G169gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(KEYINPUT62), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n853_), .ZN(G1348gat));
  NAND3_X1  g653(.A1(new_n797_), .A2(new_n677_), .A3(new_n837_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g655(.A1(new_n797_), .A2(new_n288_), .A3(new_n837_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n472_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n305_), .B2(new_n857_), .ZN(G1350gat));
  OAI211_X1 g658(.A(new_n253_), .B(new_n837_), .C1(new_n780_), .C2(new_n783_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT125), .B1(new_n860_), .B2(G190gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n797_), .A2(new_n837_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n248_), .A2(new_n310_), .ZN(new_n864_));
  OAI22_X1  g663(.A1(new_n861_), .A2(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1351gat));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n822_), .A2(new_n510_), .A3(new_n411_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n600_), .B(new_n867_), .C1(new_n780_), .C2(new_n783_), .ZN(new_n868_));
  INV_X1    g667(.A(G197gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n869_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n867_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n600_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n870_), .A2(new_n871_), .A3(new_n874_), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n677_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g676(.A(KEYINPUT63), .B(G211gat), .Z(new_n878_));
  AND3_X1   g677(.A1(new_n873_), .A2(new_n288_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n873_), .A2(new_n288_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1354gat));
  AOI21_X1  g681(.A(G218gat), .B1(new_n873_), .B2(new_n248_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n253_), .A2(G218gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT127), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n873_), .B2(new_n885_), .ZN(G1355gat));
endmodule


