//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_;
  INV_X1    g000(.A(G197gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT95), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT95), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n207_), .B2(G204gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G211gat), .A2(G218gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G211gat), .A2(G218gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT96), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT96), .ZN(new_n215_));
  INV_X1    g014(.A(new_n213_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G197gat), .A2(G204gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT95), .B(G197gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(KEYINPUT21), .B(new_n219_), .C1(new_n220_), .C2(G204gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n210_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT98), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n217_), .B(new_n214_), .C1(new_n208_), .C2(KEYINPUT97), .ZN(new_n225_));
  INV_X1    g024(.A(new_n203_), .ZN(new_n226_));
  INV_X1    g025(.A(G204gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT97), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT21), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n224_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n218_), .B1(new_n229_), .B2(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n209_), .B1(new_n208_), .B2(KEYINPUT97), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT98), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n223_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  AND2_X1   g035(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n237_), .A2(new_n238_), .B1(G141gat), .B2(G148gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT2), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(G141gat), .A3(G148gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT93), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT93), .A4(new_n247_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n250_), .A2(new_n251_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n254_), .A2(KEYINPUT1), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(new_n252_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(KEYINPUT1), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n259_), .A3(KEYINPUT91), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n258_), .B(new_n260_), .C1(KEYINPUT1), .C2(new_n254_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n240_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(new_n245_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n236_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(G228gat), .B(G233gat), .C1(new_n235_), .C2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT94), .B1(new_n255_), .B2(new_n264_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n264_), .A3(KEYINPUT94), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n236_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n225_), .A2(new_n230_), .A3(new_n224_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT98), .B1(new_n232_), .B2(new_n233_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n222_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G228gat), .A2(G233gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n266_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G78gat), .ZN(new_n277_));
  INV_X1    g076(.A(G78gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n266_), .B(new_n278_), .C1(new_n270_), .C2(new_n275_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(G106gat), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(G106gat), .B1(new_n277_), .B2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT99), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n255_), .A2(KEYINPUT94), .A3(new_n264_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n267_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n236_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT28), .B(G22gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G50gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n285_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G106gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n279_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n274_), .B(new_n273_), .C1(new_n284_), .C2(new_n236_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n278_), .B1(new_n292_), .B2(new_n266_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n277_), .A2(G106gat), .A3(new_n279_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n282_), .A2(new_n289_), .A3(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT99), .B(new_n288_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT26), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT84), .Z(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(KEYINPUT85), .A2(KEYINPUT26), .ZN(new_n306_));
  OAI21_X1  g105(.A(G190gat), .B1(KEYINPUT85), .B2(KEYINPUT26), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n304_), .B(new_n305_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT86), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT24), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT23), .B1(new_n313_), .B2(new_n302_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT87), .ZN(new_n315_));
  OR3_X1    g114(.A1(new_n313_), .A2(new_n302_), .A3(KEYINPUT23), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n317_), .B(KEYINPUT23), .C1(new_n313_), .C2(new_n302_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n310_), .A2(KEYINPUT24), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n308_), .A2(new_n312_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT88), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n314_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n313_), .A2(new_n302_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G120gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(KEYINPUT90), .ZN(new_n333_));
  INV_X1    g132(.A(G113gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(KEYINPUT90), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n331_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G113gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(G120gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n330_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT30), .B(G71gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT89), .B(G99gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT31), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n346_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n301_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n343_), .B1(new_n283_), .B2(new_n267_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT101), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n255_), .A2(new_n264_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n343_), .A2(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n343_), .B(KEYINPUT101), .C1(new_n283_), .C2(new_n267_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT4), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT103), .A3(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n362_), .A2(new_n367_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G57gat), .B(G85gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  NOR2_X1   g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT103), .ZN(new_n376_));
  INV_X1    g175(.A(new_n365_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n362_), .B2(KEYINPUT4), .ZN(new_n378_));
  INV_X1    g177(.A(new_n367_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n368_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n305_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n312_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n316_), .A2(new_n314_), .B1(new_n386_), .B2(new_n309_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n319_), .A2(new_n327_), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n385_), .A2(new_n387_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n382_), .B1(new_n235_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n273_), .A2(new_n330_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G64gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G92gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n235_), .A2(new_n392_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n235_), .A2(new_n329_), .A3(new_n321_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(KEYINPUT20), .A3(new_n397_), .A4(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT100), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n403_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n406_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n399_), .A2(new_n406_), .A3(KEYINPUT100), .A4(new_n403_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n409_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n381_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n363_), .A2(new_n379_), .A3(new_n365_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n362_), .A2(new_n367_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT33), .B1(new_n419_), .B2(new_n374_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  INV_X1    g220(.A(new_n374_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n421_), .B(new_n422_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT104), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n362_), .A2(new_n367_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n379_), .B2(new_n378_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n428_), .B2(new_n422_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n367_), .B(new_n377_), .C1(new_n362_), .C2(KEYINPUT4), .ZN(new_n430_));
  OAI211_X1 g229(.A(KEYINPUT33), .B(new_n374_), .C1(new_n430_), .C2(new_n427_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n429_), .A2(new_n415_), .A3(new_n381_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT104), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n395_), .A2(new_n397_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n404_), .A2(KEYINPUT20), .A3(new_n405_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n397_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n410_), .A2(KEYINPUT32), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n411_), .A2(new_n412_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n428_), .A2(new_n422_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n419_), .A2(new_n374_), .ZN(new_n441_));
  OAI221_X1 g240(.A(new_n438_), .B1(new_n437_), .B2(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n426_), .A2(new_n433_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n440_), .A2(new_n441_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n300_), .A2(new_n354_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n298_), .A2(new_n353_), .A3(new_n299_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n415_), .A2(KEYINPUT27), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT105), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n413_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n436_), .A2(new_n403_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n413_), .A2(new_n450_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(KEYINPUT27), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n355_), .A2(new_n443_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT64), .Z(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT65), .Z(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT6), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT7), .ZN(new_n462_));
  INV_X1    g261(.A(G99gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n290_), .A4(KEYINPUT68), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n290_), .A3(KEYINPUT68), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT7), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468_));
  XOR2_X1   g267(.A(G85gat), .B(G92gat), .Z(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT66), .B(G85gat), .ZN(new_n474_));
  INV_X1    g273(.A(G92gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n476_), .B(KEYINPUT67), .C1(new_n473_), .C2(new_n469_), .ZN(new_n477_));
  INV_X1    g276(.A(G85gat), .ZN(new_n478_));
  OR4_X1    g277(.A1(KEYINPUT67), .A2(new_n473_), .A3(new_n478_), .A4(new_n475_), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT10), .B(G99gat), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n290_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n477_), .A2(new_n479_), .A3(new_n461_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n470_), .A2(new_n471_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n472_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G64gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  XOR2_X1   g285(.A(G71gat), .B(G78gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n490_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT12), .A3(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(KEYINPUT12), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n459_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n459_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G120gat), .B(G148gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  OR2_X1    g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT71), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(KEYINPUT13), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT72), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT72), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G29gat), .B(G36gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT73), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G43gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G50gat), .ZN(new_n520_));
  INV_X1    g319(.A(G43gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n518_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G50gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526_));
  INV_X1    g325(.A(G1gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT80), .ZN(new_n535_));
  INV_X1    g334(.A(new_n525_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n532_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT81), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(KEYINPUT81), .A3(new_n537_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n515_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n525_), .B(KEYINPUT15), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n532_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n535_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n515_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(KEYINPUT82), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT82), .ZN(new_n549_));
  INV_X1    g348(.A(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n542_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n324_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n202_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n542_), .A2(new_n550_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT83), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n559_));
  NOR4_X1   g358(.A1(new_n542_), .A2(new_n550_), .A3(new_n559_), .A4(new_n554_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n555_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n456_), .A2(new_n514_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n490_), .B(new_n533_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G183gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(G211gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT78), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(KEYINPUT78), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n566_), .B(KEYINPUT75), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n573_), .B(KEYINPUT76), .ZN(new_n579_));
  OAI22_X1  g378(.A1(new_n576_), .A2(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT79), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n563_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n544_), .A2(new_n484_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n536_), .A2(new_n484_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT34), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n585_), .B(new_n586_), .C1(KEYINPUT35), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT35), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G134gat), .ZN(new_n593_));
  INV_X1    g392(.A(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT36), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n590_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n591_), .A2(new_n598_), .B1(new_n601_), .B2(new_n595_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n584_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n589_), .B(new_n590_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n599_), .A3(new_n583_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n582_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT106), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n527_), .A3(new_n445_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT38), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n599_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n582_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n444_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  OAI21_X1  g418(.A(G8gat), .B1(new_n616_), .B2(new_n455_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n455_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n528_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n619_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n620_), .B(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(KEYINPUT40), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n616_), .B2(new_n353_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n609_), .A2(G15gat), .A3(new_n353_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n615_), .B2(new_n301_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT42), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n301_), .A2(new_n634_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n609_), .B2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n581_), .A2(new_n614_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT108), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(new_n563_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G29gat), .A3(new_n444_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n456_), .B2(new_n608_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n443_), .A2(new_n355_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n447_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n353_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n455_), .B(new_n444_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n608_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(KEYINPUT43), .A3(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n514_), .A2(new_n562_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT79), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n580_), .B(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n645_), .A2(new_n652_), .A3(new_n653_), .A4(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n445_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT107), .B1(new_n658_), .B2(G29gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n643_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(G1328gat));
  XNOR2_X1  g462(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT43), .B1(new_n650_), .B2(new_n651_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n644_), .B(new_n608_), .C1(new_n646_), .C2(new_n649_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT44), .A3(new_n653_), .A4(new_n655_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n656_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n623_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT110), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n668_), .A2(new_n670_), .A3(new_n673_), .A4(new_n623_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(G36gat), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n672_), .A2(KEYINPUT111), .A3(G36gat), .A4(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n641_), .A2(new_n680_), .A3(new_n623_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n664_), .B1(new_n679_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n664_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n686_), .B(new_n683_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1329gat));
  OAI21_X1  g487(.A(new_n521_), .B1(new_n642_), .B2(new_n353_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n657_), .A2(G43gat), .A3(new_n354_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g494(.A(new_n523_), .B1(new_n657_), .B2(new_n301_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n642_), .A2(G50gat), .A3(new_n300_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT114), .ZN(G1331gat));
  INV_X1    g498(.A(new_n514_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(new_n456_), .A3(new_n561_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n581_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n651_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n445_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n613_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n445_), .A2(G57gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n705_), .B2(new_n623_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT48), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n455_), .A2(G64gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT115), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n703_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n715_), .A3(new_n354_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n705_), .A2(new_n354_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G71gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT49), .B(new_n715_), .C1(new_n705_), .C2(new_n354_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT116), .Z(G1334gat));
  AOI21_X1  g521(.A(new_n278_), .B1(new_n705_), .B2(new_n301_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n703_), .A2(new_n278_), .A3(new_n301_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n640_), .A2(new_n701_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n478_), .B1(new_n727_), .B2(new_n444_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n665_), .A2(new_n666_), .A3(new_n581_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n700_), .A2(new_n561_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n444_), .A2(new_n474_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT117), .Z(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT118), .Z(G1336gat));
  INV_X1    g534(.A(new_n727_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G92gat), .B1(new_n736_), .B2(new_n623_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n731_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n455_), .A2(new_n475_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT119), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n738_), .B2(new_n740_), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n731_), .B2(new_n353_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n480_), .A3(new_n354_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n736_), .A2(new_n290_), .A3(new_n301_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n738_), .A2(new_n301_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g552(.A1(new_n623_), .A2(new_n444_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT120), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n495_), .A2(new_n755_), .A3(KEYINPUT55), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n493_), .A2(new_n459_), .A3(new_n494_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT121), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT55), .B1(new_n495_), .B2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(KEYINPUT121), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .A4(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(KEYINPUT122), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(KEYINPUT122), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n503_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  INV_X1    g565(.A(new_n503_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n766_), .B(new_n767_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n561_), .B(new_n504_), .C1(new_n765_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n515_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n557_), .B(new_n771_), .C1(new_n770_), .C2(new_n546_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n556_), .A2(new_n557_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n559_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n556_), .A2(KEYINPUT83), .A3(new_n557_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n506_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT57), .B1(new_n778_), .B2(new_n614_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n613_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n767_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT56), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n504_), .A4(new_n776_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n776_), .B(new_n504_), .C1(new_n765_), .C2(new_n768_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(new_n651_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n581_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n562_), .A2(new_n581_), .A3(new_n511_), .A4(new_n608_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT54), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT54), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n648_), .B(new_n754_), .C1(new_n790_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797_), .B2(new_n561_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n785_), .A2(new_n788_), .A3(new_n651_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n800_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n801_), .B2(new_n581_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n648_), .A4(new_n754_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n562_), .A2(new_n334_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n798_), .B1(new_n805_), .B2(new_n806_), .ZN(G1340gat));
  INV_X1    g606(.A(KEYINPUT60), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n700_), .B2(G120gat), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n802_), .A2(new_n648_), .A3(new_n754_), .A4(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n799_), .A2(new_n804_), .A3(new_n810_), .A4(new_n514_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G120gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(KEYINPUT60), .B2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g612(.A(G127gat), .B1(new_n797_), .B2(new_n581_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n581_), .A2(G127gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n805_), .B2(new_n815_), .ZN(G1342gat));
  INV_X1    g615(.A(G134gat), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n608_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n799_), .A2(new_n804_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n796_), .B2(new_n614_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(KEYINPUT123), .A3(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1343gat));
  NOR2_X1   g624(.A1(new_n790_), .A2(new_n795_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n447_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n754_), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n828_), .A2(G141gat), .A3(new_n562_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G141gat), .B1(new_n828_), .B2(new_n562_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1344gat));
  OR3_X1    g630(.A1(new_n828_), .A2(G148gat), .A3(new_n700_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G148gat), .B1(new_n828_), .B2(new_n700_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1345gat));
  NAND3_X1  g633(.A1(new_n827_), .A2(new_n581_), .A3(new_n754_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  NOR3_X1   g636(.A1(new_n828_), .A2(new_n594_), .A3(new_n608_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n828_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n613_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n594_), .B2(new_n840_), .ZN(G1347gat));
  NOR2_X1   g640(.A1(new_n826_), .A2(new_n446_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n455_), .A2(new_n445_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n561_), .A3(new_n389_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n561_), .A2(new_n843_), .A3(new_n354_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT124), .Z(new_n848_));
  OAI211_X1 g647(.A(new_n300_), .B(new_n848_), .C1(new_n790_), .C2(new_n795_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT125), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n802_), .A2(new_n851_), .A3(new_n300_), .A4(new_n848_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(G169gat), .A3(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(KEYINPUT62), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(KEYINPUT62), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n846_), .B1(new_n854_), .B2(new_n855_), .ZN(G1348gat));
  NAND3_X1  g655(.A1(new_n842_), .A2(new_n514_), .A3(new_n843_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n313_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n845_), .A2(new_n305_), .A3(new_n581_), .A4(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n844_), .A2(new_n655_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n859_), .A2(G183gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(G1350gat));
  OAI21_X1  g663(.A(G190gat), .B1(new_n844_), .B2(new_n608_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n613_), .A2(new_n383_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n844_), .B2(new_n866_), .ZN(G1351gat));
  NAND3_X1  g666(.A1(new_n827_), .A2(new_n561_), .A3(new_n843_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n827_), .A2(new_n843_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n227_), .A3(new_n514_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G204gat), .B1(new_n870_), .B2(new_n700_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1353gat));
  NAND3_X1  g673(.A1(new_n827_), .A2(new_n581_), .A3(new_n843_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT63), .B(G211gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n875_), .B2(new_n878_), .ZN(G1354gat));
  XOR2_X1   g678(.A(KEYINPUT127), .B(G218gat), .Z(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n870_), .A2(new_n608_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n871_), .A2(new_n613_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1355gat));
endmodule


