//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  INV_X1    g014(.A(new_n206_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n209_), .A2(KEYINPUT66), .A3(new_n206_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n205_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n211_), .B1(new_n221_), .B2(KEYINPUT67), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n223_), .A3(new_n212_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n205_), .B1(G106gat), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G85gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G92gat), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n230_), .A2(new_n231_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n234_), .B(KEYINPUT65), .Z(new_n235_));
  AOI21_X1  g034(.A(new_n227_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n225_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  INV_X1    g037(.A(new_n236_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n220_), .A2(new_n223_), .A3(new_n212_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n223_), .B1(new_n220_), .B2(new_n212_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n211_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n238_), .B(new_n239_), .C1(new_n242_), .C2(new_n214_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT69), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n203_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n237_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n257_), .B(new_n214_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT70), .B1(new_n260_), .B2(new_n213_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n239_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n250_), .A2(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n256_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n254_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n251_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n203_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G120gat), .B(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT5), .B(G176gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n265_), .A2(new_n268_), .A3(KEYINPUT71), .A4(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n265_), .A2(new_n268_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT13), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n282_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT72), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT85), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n291_), .A2(new_n297_), .A3(KEYINPUT1), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(G141gat), .ZN(new_n301_));
  INV_X1    g100(.A(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT86), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(KEYINPUT3), .ZN(new_n307_));
  OR3_X1    g106(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n292_), .A2(new_n295_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT87), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n306_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(KEYINPUT91), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n316_), .A2(new_n320_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n325_), .B2(KEYINPUT4), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n327_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(new_n232_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n329_), .A2(KEYINPUT33), .A3(new_n335_), .A4(new_n330_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(KEYINPUT92), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(new_n231_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT18), .B(G64gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT23), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT82), .Z(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n349_), .B2(KEYINPUT24), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT83), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT83), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT24), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT81), .Z(new_n358_));
  NAND4_X1  g157(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .A4(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n347_), .B1(G183gat), .B2(G190gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  INV_X1    g160(.A(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n363_), .A3(new_n353_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT88), .B(G197gat), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n366_), .A2(G204gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(G197gat), .B2(G204gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G211gat), .B(G218gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n270_), .A2(G197gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n366_), .B2(new_n270_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n370_), .B(new_n371_), .C1(KEYINPUT21), .C2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n371_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(KEYINPUT21), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n365_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n353_), .A2(KEYINPUT24), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT90), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(KEYINPUT90), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n349_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n347_), .B(new_n357_), .C1(new_n349_), .C2(KEYINPUT24), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n364_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(KEYINPUT20), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n377_), .A2(new_n385_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT20), .B(new_n392_), .C1(new_n365_), .C2(new_n378_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(new_n389_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n345_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n345_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n390_), .B(new_n396_), .C1(new_n389_), .C2(new_n393_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n326_), .A2(new_n327_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n335_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .A4(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n391_), .A2(new_n394_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n389_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n389_), .B2(new_n387_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n406_), .B2(new_n403_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n336_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n331_), .A2(new_n335_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n402_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n365_), .B(KEYINPUT30), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G71gat), .B(G99gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n319_), .B(KEYINPUT31), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n412_), .A2(new_n413_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n414_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n420_), .B(new_n421_), .C1(new_n423_), .C2(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n419_), .B1(new_n422_), .B2(new_n414_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n420_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n431_));
  XOR2_X1   g230(.A(G22gat), .B(G50gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT28), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n431_), .B(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n378_), .B1(new_n316_), .B2(KEYINPUT29), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G78gat), .B(G106gat), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n434_), .B1(new_n440_), .B2(KEYINPUT89), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n437_), .B(new_n439_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n430_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n409_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n336_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n345_), .B(KEYINPUT93), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n406_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n397_), .A3(KEYINPUT27), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n398_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n448_), .A2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n443_), .A2(new_n444_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n430_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n429_), .A2(new_n445_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n411_), .A2(new_n446_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(G197gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT79), .B(G169gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n468_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n475_));
  XOR2_X1   g274(.A(G1gat), .B(G8gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT76), .ZN(new_n477_));
  INV_X1    g276(.A(G15gat), .ZN(new_n478_));
  INV_X1    g277(.A(G22gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G15gat), .A2(G22gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G1gat), .A2(G8gat), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n480_), .A2(new_n481_), .B1(KEYINPUT14), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n477_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n475_), .A2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n477_), .A2(new_n483_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n477_), .A2(new_n483_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n474_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n474_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT80), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n467_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n467_), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT80), .B(new_n501_), .C1(new_n492_), .C2(new_n497_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n290_), .A2(new_n463_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n262_), .A2(new_n475_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n244_), .A2(new_n474_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT35), .A3(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n505_), .A2(new_n506_), .A3(new_n512_), .A4(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G190gat), .B(G218gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G134gat), .B(G162gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT74), .Z(new_n520_));
  NOR2_X1   g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n517_), .B(KEYINPUT36), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n514_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT75), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT75), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n514_), .B2(new_n523_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT96), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT97), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(G211gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT16), .B(G183gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT69), .B1(new_n534_), .B2(KEYINPUT17), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT77), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n250_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n536_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n488_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n540_), .B1(KEYINPUT17), .B2(new_n534_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n488_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n530_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n504_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n202_), .B1(new_n546_), .B2(new_n448_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n528_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n522_), .A2(KEYINPUT37), .A3(new_n524_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n543_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n463_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n289_), .B(KEYINPUT73), .ZN(new_n558_));
  INV_X1    g357(.A(new_n503_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n448_), .A2(new_n202_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n547_), .B1(new_n564_), .B2(KEYINPUT38), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(KEYINPUT38), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n564_), .A2(KEYINPUT98), .A3(KEYINPUT38), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(G1324gat));
  NAND2_X1  g369(.A1(new_n546_), .A2(new_n457_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(G8gat), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n457_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n562_), .A2(G8gat), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n574_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(G1325gat));
  AOI21_X1  g380(.A(new_n478_), .B1(new_n546_), .B2(new_n430_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT41), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n430_), .A2(new_n478_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n585_), .C1(new_n560_), .C2(new_n586_), .ZN(G1326gat));
  OAI21_X1  g386(.A(G22gat), .B1(new_n545_), .B2(new_n459_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT42), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n445_), .A2(new_n479_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT100), .Z(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n560_), .B2(new_n591_), .ZN(G1327gat));
  INV_X1    g391(.A(KEYINPUT102), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n289_), .A2(new_n543_), .A3(new_n559_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT101), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT43), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n411_), .A2(new_n446_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n458_), .A2(new_n462_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n597_), .B(new_n551_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n552_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(KEYINPUT101), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT44), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n596_), .A2(new_n602_), .A3(KEYINPUT44), .A4(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n448_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n593_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n606_), .A2(KEYINPUT102), .A3(new_n448_), .A4(new_n607_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(G29gat), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n529_), .A2(new_n553_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n504_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(G29gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT103), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT104), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1328gat));
  OAI21_X1  g422(.A(G36gat), .B1(new_n608_), .B2(new_n575_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n614_), .A2(G36gat), .A3(new_n575_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT45), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT46), .Z(G1329gat));
  NOR3_X1   g428(.A1(new_n614_), .A2(G43gat), .A3(new_n429_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n606_), .A2(new_n430_), .A3(new_n607_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(G43gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g432(.A(G50gat), .B1(new_n608_), .B2(new_n459_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n614_), .A2(G50gat), .A3(new_n459_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1331gat));
  NOR3_X1   g435(.A1(new_n558_), .A2(new_n463_), .A3(new_n559_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n544_), .ZN(new_n638_));
  INV_X1    g437(.A(G57gat), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n609_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n290_), .A2(new_n503_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n557_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n448_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n640_), .B1(new_n647_), .B2(new_n639_), .ZN(G1332gat));
  OAI21_X1  g447(.A(G64gat), .B1(new_n638_), .B2(new_n575_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT48), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n575_), .A2(G64gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n643_), .B2(new_n651_), .ZN(G1333gat));
  OAI21_X1  g451(.A(G71gat), .B1(new_n638_), .B2(new_n429_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT49), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n429_), .A2(G71gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT106), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n644_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(KEYINPUT107), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1334gat));
  OAI21_X1  g461(.A(G78gat), .B1(new_n638_), .B2(new_n459_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT50), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n459_), .A2(G78gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n643_), .B2(new_n665_), .ZN(G1335gat));
  NAND2_X1  g465(.A1(new_n637_), .A2(new_n613_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n232_), .B1(new_n667_), .B2(new_n609_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n553_), .B(new_n641_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n609_), .A2(new_n228_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT108), .ZN(G1336gat));
  NAND3_X1  g472(.A1(new_n637_), .A2(new_n457_), .A3(new_n613_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n457_), .A2(G92gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT109), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n674_), .A2(new_n231_), .B1(new_n669_), .B2(new_n676_), .ZN(G1337gat));
  NOR3_X1   g476(.A1(new_n667_), .A2(new_n226_), .A3(new_n429_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n430_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G99gat), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g480(.A1(new_n667_), .A2(G106gat), .A3(new_n459_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n669_), .A2(new_n445_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT52), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G106gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G106gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g487(.A1(new_n283_), .A2(new_n503_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n554_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n554_), .B2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n278_), .B2(new_n559_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT111), .B(new_n503_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n254_), .A2(new_n255_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(KEYINPUT55), .A3(new_n253_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n244_), .A2(new_n252_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n256_), .A2(new_n703_), .A3(new_n264_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n203_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT55), .B1(new_n701_), .B2(new_n253_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(new_n705_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n280_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT56), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n699_), .B(new_n700_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n490_), .A2(new_n491_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n495_), .A2(new_n496_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n467_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n498_), .B2(new_n467_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n282_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n705_), .A2(new_n702_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n707_), .B1(new_n265_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n706_), .A2(new_n707_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n273_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT56), .B1(new_n728_), .B2(KEYINPUT113), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n700_), .B1(new_n731_), .B2(new_n699_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n529_), .B1(new_n722_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT57), .B(new_n529_), .C1(new_n722_), .C2(new_n732_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT118), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT117), .B1(new_n728_), .B2(KEYINPUT56), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT56), .B(new_n280_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n710_), .A2(new_n742_), .A3(new_n712_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n278_), .A2(new_n720_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT58), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n739_), .B1(new_n747_), .B2(new_n552_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n743_), .A2(new_n741_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n745_), .B1(new_n749_), .B2(new_n740_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT118), .B(new_n551_), .C1(new_n750_), .C2(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT58), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n733_), .A2(KEYINPUT116), .A3(new_n734_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n737_), .A2(new_n738_), .A3(new_n753_), .A4(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n695_), .B1(new_n755_), .B2(new_n543_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n609_), .A2(new_n457_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n460_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT119), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n733_), .A2(KEYINPUT116), .A3(new_n734_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT116), .B1(new_n733_), .B2(new_n734_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n753_), .A2(new_n738_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n553_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n762_), .B(new_n759_), .C1(new_n767_), .C2(new_n695_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n761_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G113gat), .B1(new_n769_), .B2(new_n559_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n755_), .A2(new_n543_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n760_), .B1(new_n771_), .B2(new_n694_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n753_), .A2(new_n738_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n735_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n543_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n694_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n760_), .A2(KEYINPUT59), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n773_), .A2(KEYINPUT59), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n559_), .A2(G113gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n779_), .B2(new_n780_), .ZN(G1340gat));
  NOR2_X1   g580(.A1(new_n289_), .A2(KEYINPUT60), .ZN(new_n782_));
  MUX2_X1   g581(.A(new_n782_), .B(KEYINPUT60), .S(G120gat), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n769_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n773_), .A2(KEYINPUT59), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  INV_X1    g585(.A(new_n558_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n777_), .A2(new_n778_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G120gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n779_), .B2(new_n787_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n790_), .B2(new_n791_), .ZN(G1341gat));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n553_), .B(new_n788_), .C1(new_n772_), .C2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G127gat), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n543_), .A2(G127gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n769_), .A2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1342gat));
  NAND2_X1  g600(.A1(new_n769_), .A2(new_n530_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n803_));
  INV_X1    g602(.A(G134gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n779_), .A2(G134gat), .A3(new_n551_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n530_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n761_), .B2(new_n768_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT122), .B1(new_n808_), .B2(G134gat), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n809_), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n756_), .A2(new_n461_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n757_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n503_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(new_n301_), .ZN(G1344gat));
  NOR2_X1   g613(.A1(new_n812_), .A2(new_n558_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n302_), .ZN(G1345gat));
  OAI21_X1  g615(.A(KEYINPUT123), .B1(new_n812_), .B2(new_n543_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n811_), .A2(new_n818_), .A3(new_n553_), .A4(new_n757_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1346gat));
  NAND2_X1  g622(.A1(new_n551_), .A2(G162gat), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n756_), .A2(new_n461_), .A3(new_n807_), .A4(new_n758_), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n812_), .A2(new_n824_), .B1(new_n825_), .B2(G162gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT124), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n448_), .A2(new_n575_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n460_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n777_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G169gat), .B1(new_n831_), .B2(new_n503_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT62), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n559_), .A2(new_n361_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT125), .Z(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n831_), .B2(new_n835_), .ZN(G1348gat));
  INV_X1    g635(.A(new_n831_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G176gat), .B1(new_n837_), .B2(new_n290_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n756_), .A2(new_n445_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n558_), .A2(new_n362_), .A3(new_n429_), .A4(new_n829_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  NOR3_X1   g640(.A1(new_n831_), .A2(new_n543_), .A3(new_n355_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n839_), .A2(new_n553_), .A3(new_n430_), .A4(new_n828_), .ZN(new_n843_));
  INV_X1    g642(.A(G183gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(G1350gat));
  OAI21_X1  g644(.A(G190gat), .B1(new_n831_), .B2(new_n552_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n530_), .A2(new_n356_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT126), .Z(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n831_), .B2(new_n848_), .ZN(G1351gat));
  NOR3_X1   g648(.A1(new_n756_), .A2(new_n461_), .A3(new_n829_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n559_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n787_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g653(.A1(new_n850_), .A2(new_n553_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n855_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT63), .B(G211gat), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n855_), .B2(new_n857_), .ZN(G1354gat));
  XNOR2_X1  g657(.A(KEYINPUT127), .B(G218gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n850_), .B2(new_n530_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n551_), .A2(new_n859_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n850_), .B2(new_n861_), .ZN(G1355gat));
endmodule


