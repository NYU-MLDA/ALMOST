//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT22), .B(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(new_n210_), .C1(G183gat), .C2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n206_), .B(new_n211_), .C1(new_n212_), .C2(new_n205_), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G190gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT91), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT91), .B1(new_n215_), .B2(new_n217_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT25), .B(G183gat), .Z(new_n220_));
  NOR3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n212_), .A3(new_n205_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n213_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G197gat), .A2(G204gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT21), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233_));
  INV_X1    g032(.A(new_n231_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n229_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n234_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n236_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT87), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n232_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n237_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n203_), .B1(new_n228_), .B2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n224_), .A2(new_n226_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n215_), .A2(new_n217_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT81), .B1(new_n220_), .B2(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n215_), .A2(new_n217_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT25), .B(G183gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT87), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n241_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n255_), .A3(new_n237_), .A4(new_n213_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT19), .Z(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT90), .Z(new_n260_));
  OR2_X1    g059(.A1(new_n228_), .A2(new_n243_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(KEYINPUT20), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n213_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n243_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n257_), .A2(new_n260_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n202_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n257_), .A2(new_n260_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n263_), .B2(new_n243_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n259_), .B1(new_n261_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n270_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n260_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n244_), .B2(new_n256_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n261_), .A2(new_n264_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n271_), .A3(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n261_), .A2(new_n264_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n270_), .B1(new_n285_), .B2(new_n281_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT27), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT100), .B1(new_n279_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n286_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n289_), .A2(new_n202_), .B1(new_n272_), .B2(new_n278_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT100), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT82), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n263_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n252_), .A2(KEYINPUT30), .A3(new_n213_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G227gat), .ZN(new_n303_));
  INV_X1    g102(.A(G233gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n302_), .A2(new_n305_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n298_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G134gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G127gat), .ZN(new_n313_));
  INV_X1    g112(.A(G127gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G134gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n311_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT83), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n310_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT31), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT84), .ZN(new_n326_));
  INV_X1    g125(.A(new_n302_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n305_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n306_), .A3(new_n297_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n309_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n325_), .B(KEYINPUT84), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n309_), .B2(new_n330_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT0), .ZN(new_n337_));
  INV_X1    g136(.A(G57gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G85gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344_));
  INV_X1    g143(.A(G141gat), .ZN(new_n345_));
  INV_X1    g144(.A(G148gat), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .A4(KEYINPUT85), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n350_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G155gat), .B(G162gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G141gat), .B(G148gat), .Z(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n357_), .B(new_n358_), .C1(KEYINPUT1), .C2(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n324_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n343_), .B1(new_n361_), .B2(KEYINPUT4), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n356_), .A2(new_n319_), .A3(new_n323_), .A4(new_n359_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n324_), .A2(new_n360_), .A3(KEYINPUT93), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n367_), .B2(KEYINPUT4), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n343_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n341_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT98), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT98), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(new_n341_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n342_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n339_), .B(G85gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n374_), .B(new_n375_), .C1(new_n377_), .C2(new_n362_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n373_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT86), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n243_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT88), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n243_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G228gat), .A3(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n380_), .A2(new_n387_), .A3(new_n243_), .A4(new_n382_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n384_), .A2(new_n386_), .A3(new_n392_), .A4(new_n388_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT28), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(new_n396_), .ZN(new_n397_));
  AND4_X1   g196(.A1(KEYINPUT89), .A2(new_n391_), .A3(new_n393_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n400_), .A2(new_n397_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NOR4_X1   g201(.A1(new_n293_), .A2(new_n335_), .A3(new_n379_), .A4(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n368_), .A2(new_n369_), .A3(new_n341_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(KEYINPUT98), .B2(new_n370_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n290_), .A2(new_n405_), .A3(new_n373_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n334_), .B1(new_n406_), .B2(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n378_), .A2(KEYINPUT95), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n367_), .A2(KEYINPUT4), .ZN(new_n409_));
  INV_X1    g208(.A(new_n362_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n374_), .A4(new_n375_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n404_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n378_), .B2(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n367_), .A2(new_n343_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n342_), .B1(new_n361_), .B2(KEYINPUT4), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n419_), .B(new_n341_), .C1(new_n377_), .C2(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n421_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .A4(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n265_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT96), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n265_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n273_), .A2(new_n277_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n426_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n379_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n398_), .A2(new_n401_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n423_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n407_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT99), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n407_), .A2(new_n434_), .A3(KEYINPUT99), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n403_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G134gat), .B(G162gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT72), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G190gat), .ZN(new_n442_));
  INV_X1    g241(.A(G218gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT36), .ZN(new_n445_));
  INV_X1    g244(.A(G50gat), .ZN(new_n446_));
  INV_X1    g245(.A(G43gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448_));
  INV_X1    g247(.A(G36gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G29gat), .ZN(new_n450_));
  INV_X1    g249(.A(G29gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G36gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n452_), .A3(new_n448_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n447_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n450_), .A2(new_n452_), .A3(new_n448_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n457_), .A2(new_n453_), .A3(G43gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n446_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n455_), .A3(new_n447_), .ZN(new_n460_));
  OAI21_X1  g259(.A(G43gat), .B1(new_n457_), .B2(new_n453_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(G50gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT10), .B(G99gat), .Z(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G85gat), .B(G92gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT9), .ZN(new_n468_));
  INV_X1    g267(.A(G92gat), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n340_), .A2(new_n469_), .A3(KEYINPUT9), .ZN(new_n470_));
  AND3_X1   g269(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n473_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT8), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n467_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT64), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT64), .B1(new_n471_), .B2(new_n472_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(new_n489_), .B2(new_n467_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n481_), .B1(new_n490_), .B2(KEYINPUT65), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT65), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n492_), .B(new_n480_), .C1(new_n489_), .C2(new_n467_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n463_), .B(new_n474_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n474_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n481_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n467_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n498_), .B2(new_n492_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n493_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n460_), .A2(new_n461_), .A3(G50gat), .ZN(new_n503_));
  AOI21_X1  g302(.A(G50gat), .B1(new_n460_), .B2(new_n461_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n459_), .A2(KEYINPUT15), .A3(new_n462_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n494_), .B1(new_n501_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n511_), .B(KEYINPUT34), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n508_), .A2(KEYINPUT71), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n508_), .B2(KEYINPUT71), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n512_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(KEYINPUT71), .A3(new_n513_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT35), .A3(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n444_), .A2(KEYINPUT36), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n516_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n445_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n439_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G176gat), .B(G204gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G64gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G57gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(G57gat), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n338_), .A2(G64gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT11), .B1(new_n533_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G71gat), .B(G78gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT66), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n540_), .A2(KEYINPUT66), .A3(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n538_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OR3_X1    g344(.A1(new_n540_), .A2(KEYINPUT66), .A3(new_n541_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n474_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n474_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  INV_X1    g352(.A(new_n548_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n550_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n501_), .A2(new_n548_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n549_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n531_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n561_), .A3(new_n531_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(KEYINPUT68), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  INV_X1    g365(.A(new_n564_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n562_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n568_), .A3(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT76), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(KEYINPUT17), .B2(new_n580_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583_));
  INV_X1    g382(.A(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT14), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G1gat), .B(G8gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n548_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n581_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT77), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT77), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G169gat), .ZN(new_n603_));
  INV_X1    g402(.A(G197gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n507_), .A2(new_n589_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n463_), .A2(new_n589_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n463_), .A2(new_n589_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT80), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n606_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(KEYINPUT80), .B(new_n605_), .C1(new_n611_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n574_), .A2(new_n601_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n525_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n379_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n516_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT73), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n524_), .B(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n597_), .A2(KEYINPUT78), .A3(new_n599_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT78), .B1(new_n597_), .B2(new_n599_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n629_), .A2(KEYINPUT79), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT79), .B1(new_n629_), .B2(new_n633_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n573_), .B(KEYINPUT69), .Z(new_n637_));
  INV_X1    g436(.A(new_n293_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n335_), .A2(new_n379_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n433_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n407_), .A2(new_n434_), .A3(KEYINPUT99), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT99), .B1(new_n407_), .B2(new_n434_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n618_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n637_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n636_), .A2(new_n584_), .A3(new_n379_), .A4(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT101), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n624_), .B1(new_n649_), .B2(new_n650_), .ZN(G1324gat));
  OAI21_X1  g450(.A(G8gat), .B1(new_n620_), .B2(new_n638_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT39), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n636_), .A2(new_n646_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n293_), .A2(new_n585_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n622_), .A2(new_n335_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(G15gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(G15gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n659_), .A2(G15gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT103), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT41), .A3(new_n661_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n654_), .A2(G15gat), .A3(new_n335_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n667_), .A3(new_n668_), .ZN(G1326gat));
  OAI21_X1  g468(.A(G22gat), .B1(new_n622_), .B2(new_n433_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n433_), .A2(G22gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n654_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n633_), .A2(new_n674_), .A3(new_n524_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n524_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT104), .B1(new_n632_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(new_n643_), .A3(new_n644_), .A4(new_n573_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n379_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n633_), .A2(new_n573_), .A3(new_n644_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT37), .B1(new_n522_), .B2(KEYINPUT73), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n524_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n516_), .A2(new_n520_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n521_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n626_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n628_), .A3(new_n445_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n439_), .A2(KEYINPUT43), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n643_), .B2(new_n629_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n683_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(new_n451_), .A3(new_n623_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n683_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n681_), .B1(new_n697_), .B2(new_n700_), .ZN(G1328gat));
  NAND2_X1  g500(.A1(new_n695_), .A2(new_n293_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n691_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n643_), .A2(new_n629_), .A3(new_n693_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n682_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(KEYINPUT44), .ZN(new_n706_));
  OAI21_X1  g505(.A(G36gat), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n638_), .A2(G36gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT45), .B1(new_n679_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n645_), .A2(new_n574_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n678_), .A4(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n707_), .A2(KEYINPUT46), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT107), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n707_), .A2(new_n714_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT46), .B1(new_n718_), .B2(KEYINPUT105), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n707_), .A2(new_n720_), .A3(new_n714_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n638_), .B1(new_n705_), .B2(KEYINPUT44), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n449_), .B1(new_n723_), .B2(new_n700_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n710_), .A2(new_n713_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT105), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  AND4_X1   g526(.A1(new_n717_), .A2(new_n726_), .A3(new_n727_), .A4(new_n721_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n716_), .B1(new_n722_), .B2(new_n728_), .ZN(G1329gat));
  OAI21_X1  g528(.A(new_n447_), .B1(new_n679_), .B2(new_n335_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n695_), .A2(G43gat), .A3(new_n334_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n706_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n680_), .B2(new_n402_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n696_), .A2(new_n446_), .A3(new_n433_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n700_), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n637_), .A2(new_n525_), .A3(new_n618_), .A4(new_n632_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT111), .B(G57gat), .Z(new_n738_));
  OR3_X1    g537(.A1(new_n737_), .A2(new_n623_), .A3(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n634_), .A2(new_n574_), .A3(new_n635_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n634_), .A2(KEYINPUT108), .A3(new_n574_), .A4(new_n635_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n643_), .A2(new_n618_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT109), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n742_), .A2(new_n379_), .A3(new_n743_), .A4(new_n745_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT110), .A3(new_n338_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT110), .B1(new_n746_), .B2(new_n338_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n739_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT112), .B(new_n739_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1332gat));
  OAI21_X1  g552(.A(G64gat), .B1(new_n737_), .B2(new_n638_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT48), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n293_), .A2(new_n532_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n737_), .B2(new_n335_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n335_), .A2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n756_), .B2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n737_), .B2(new_n433_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n433_), .A2(G78gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n756_), .B2(new_n767_), .ZN(G1335gat));
  AND2_X1   g567(.A1(new_n637_), .A2(new_n678_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n745_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n340_), .A3(new_n379_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n692_), .A2(new_n694_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n574_), .A2(new_n618_), .A3(new_n633_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n623_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n777_), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n469_), .A3(new_n293_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G92gat), .B1(new_n776_), .B2(new_n638_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n776_), .B2(new_n335_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n334_), .A2(new_n464_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n770_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n465_), .A3(new_n402_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n775_), .A2(new_n402_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G106gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT52), .B(new_n465_), .C1(new_n775_), .C2(new_n402_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR4_X1   g591(.A1(new_n293_), .A2(new_n335_), .A3(new_n623_), .A4(new_n402_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n524_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n616_), .A2(new_n617_), .A3(new_n564_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n549_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n558_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n557_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n551_), .B(KEYINPUT55), .C1(new_n555_), .C2(new_n556_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n530_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n531_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n807_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n801_), .A2(new_n557_), .B1(new_n799_), .B2(new_n558_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n803_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT114), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n798_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n609_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n608_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n607_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n606_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n614_), .B2(new_n606_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n565_), .A2(new_n568_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n797_), .B1(new_n814_), .B2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n820_), .A2(new_n564_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n805_), .B2(new_n812_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n824_), .B(KEYINPUT58), .C1(new_n805_), .C2(new_n812_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n685_), .A2(new_n827_), .A3(new_n690_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n804_), .A2(KEYINPUT114), .A3(new_n807_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n832_), .B2(new_n798_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n833_), .B2(new_n676_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n633_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n691_), .A2(new_n618_), .A3(new_n573_), .A4(new_n632_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n574_), .A2(new_n644_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n632_), .A4(new_n691_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n835_), .A2(new_n836_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT117), .B(new_n633_), .C1(new_n830_), .C2(new_n834_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n795_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n805_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n808_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n813_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n798_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n822_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n796_), .B1(new_n851_), .B2(new_n524_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT115), .A3(new_n823_), .A4(new_n829_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n601_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n841_), .A2(new_n838_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n793_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n844_), .B1(new_n857_), .B2(KEYINPUT59), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n618_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n618_), .A2(G113gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n857_), .B2(new_n861_), .ZN(G1340gat));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n858_), .B2(new_n637_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n857_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(KEYINPUT60), .B2(new_n864_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n867_), .A2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n866_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n863_), .B1(new_n865_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n856_), .B2(new_n793_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n637_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n844_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n873_), .B(KEYINPUT119), .C1(new_n879_), .C2(new_n864_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n880_), .ZN(G1341gat));
  OAI21_X1  g680(.A(G127gat), .B1(new_n859_), .B2(new_n601_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n866_), .A2(new_n314_), .A3(new_n632_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1342gat));
  OAI21_X1  g683(.A(G134gat), .B1(new_n859_), .B2(new_n691_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n866_), .A2(new_n312_), .A3(new_n524_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1343gat));
  NAND2_X1  g686(.A1(new_n335_), .A2(new_n402_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n888_), .A2(new_n293_), .A3(new_n623_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n856_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n618_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT120), .B(G141gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT121), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n891_), .B(new_n893_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n878_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n346_), .ZN(G1345gat));
  NAND3_X1  g695(.A1(new_n856_), .A2(new_n632_), .A3(new_n889_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT122), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(KEYINPUT122), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n900_), .B(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n890_), .B2(new_n676_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT123), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n890_), .A2(new_n904_), .A3(new_n691_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1347gat));
  NAND2_X1  g707(.A1(new_n842_), .A2(new_n843_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n639_), .A2(new_n293_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n402_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n910_), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n204_), .A3(new_n644_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n909_), .A2(new_n644_), .A3(new_n912_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n918_), .A2(new_n919_), .A3(G169gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n918_), .B2(G169gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n917_), .B1(new_n920_), .B2(new_n921_), .ZN(G1348gat));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n574_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n402_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n878_), .A2(new_n205_), .A3(new_n911_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n923_), .A2(new_n205_), .B1(new_n924_), .B2(new_n925_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n633_), .A2(new_n911_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G183gat), .B1(new_n924_), .B2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n601_), .A2(new_n250_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n916_), .B2(new_n929_), .ZN(G1350gat));
  INV_X1    g729(.A(new_n915_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n913_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G190gat), .B1(new_n932_), .B2(new_n691_), .ZN(new_n933_));
  OR3_X1    g732(.A1(new_n676_), .A2(new_n219_), .A3(new_n218_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n932_), .B2(new_n934_), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n888_), .A2(new_n379_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n293_), .B1(new_n936_), .B2(KEYINPUT125), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(KEYINPUT125), .B2(new_n936_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n856_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT126), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n856_), .A2(new_n941_), .A3(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n644_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT127), .B(G197gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1352gat));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n637_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g747(.A(new_n601_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n943_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n950_), .B(new_n952_), .ZN(G1354gat));
  NAND3_X1  g752(.A1(new_n943_), .A2(new_n443_), .A3(new_n524_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n691_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n443_), .ZN(G1355gat));
endmodule


