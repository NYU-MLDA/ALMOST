//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT8), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n205_), .B(new_n206_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n216_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n210_), .B1(new_n221_), .B2(KEYINPUT66), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n215_), .A2(new_n223_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(new_n206_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n212_), .A2(new_n214_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n216_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n222_), .A2(new_n224_), .B1(KEYINPUT8), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT65), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  AND2_X1   g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(new_n231_), .ZN(new_n237_));
  AOI21_X1  g036(.A(G106gat), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n205_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n215_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n230_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT66), .B1(new_n227_), .B2(new_n228_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n210_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n224_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n229_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n242_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G29gat), .B(G36gat), .Z(new_n251_));
  XOR2_X1   g050(.A(G43gat), .B(G50gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G29gat), .B(G36gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n243_), .A2(new_n250_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n230_), .B2(new_n242_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n248_), .A2(KEYINPUT71), .A3(new_n249_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT77), .B(KEYINPUT15), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n257_), .B(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT35), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT76), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT76), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n258_), .A2(new_n264_), .A3(new_n272_), .A4(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n267_), .A2(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G190gat), .B(G218gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(KEYINPUT36), .A3(new_n278_), .A4(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(KEYINPUT36), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n271_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n275_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n283_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n282_), .B1(new_n286_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT37), .ZN(new_n292_));
  XOR2_X1   g091(.A(G127gat), .B(G155gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G183gat), .B(G211gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT80), .B1(new_n297_), .B2(KEYINPUT17), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n298_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT69), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT11), .ZN(new_n311_));
  XOR2_X1   g110(.A(G71gat), .B(G78gat), .Z(new_n312_));
  NOR3_X1   g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n310_), .A2(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n312_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n311_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n308_), .A2(new_n318_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT37), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n282_), .B(new_n323_), .C1(new_n286_), .C2(new_n290_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n292_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n309_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT11), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n317_), .A3(new_n312_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n314_), .A2(new_n315_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n243_), .A2(new_n331_), .A3(new_n250_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G230gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT64), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n202_), .B(new_n242_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT68), .B1(new_n248_), .B2(new_n249_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n318_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT12), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n318_), .A2(KEYINPUT12), .A3(new_n260_), .A4(new_n261_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n318_), .B(KEYINPUT70), .C1(new_n337_), .C2(new_n338_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n331_), .B1(new_n243_), .B2(new_n250_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n334_), .B(new_n344_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G120gat), .B(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT5), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G176gat), .B(G204gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n343_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT72), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n343_), .A2(new_n348_), .A3(new_n356_), .A4(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT73), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n362_), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n366_));
  OR2_X1    g165(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT73), .B(new_n359_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n366_), .B(new_n367_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n325_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT81), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(KEYINPUT81), .ZN(new_n375_));
  INV_X1    g174(.A(new_n305_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n257_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n305_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G229gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n263_), .A2(new_n305_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n377_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n384_), .B2(new_n381_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G141gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G169gat), .B(G197gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT82), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n385_), .A2(KEYINPUT82), .A3(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT23), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(G183gat), .B2(G190gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G169gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT25), .B(G183gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(G190gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n405_), .A2(new_n406_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(KEYINPUT23), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT91), .ZN(new_n415_));
  OR3_X1    g214(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n410_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT92), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT92), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n410_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n404_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(G197gat), .A2(G204gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G197gat), .A2(G204gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(KEYINPUT21), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G211gat), .B(G218gat), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT21), .B1(new_n424_), .B2(new_n425_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n426_), .B(new_n427_), .C1(new_n429_), .C2(KEYINPUT89), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n425_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT21), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT89), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n428_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n423_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n414_), .A2(new_n416_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n409_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n441_), .A2(new_n407_), .A3(KEYINPUT85), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT26), .ZN(new_n444_));
  INV_X1    g243(.A(G190gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT83), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G190gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT84), .B(new_n405_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n450_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(G190gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n444_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT84), .B1(new_n455_), .B2(new_n405_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n443_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G183gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n399_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n402_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n436_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT20), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n397_), .B1(new_n437_), .B2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G8gat), .B(G36gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT18), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n457_), .A2(new_n461_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n435_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n423_), .A2(new_n436_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n397_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n464_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT27), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n435_), .A2(KEYINPUT90), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(new_n428_), .C1(new_n430_), .C2(new_n434_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n403_), .A3(new_n419_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n471_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n397_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n438_), .A2(KEYINPUT91), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n421_), .B1(new_n486_), .B2(new_n410_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n422_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n403_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n435_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n405_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n451_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n494_), .A2(new_n443_), .B1(new_n402_), .B2(new_n460_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n469_), .B1(new_n495_), .B2(new_n436_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(new_n496_), .A3(new_n473_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n483_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n468_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n476_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT27), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n464_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n468_), .B1(new_n464_), .B2(new_n474_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT98), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n473_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT20), .B(new_n473_), .C1(new_n495_), .C2(new_n436_), .ZN(new_n507_));
  AOI211_X1 g306(.A(new_n435_), .B(new_n404_), .C1(new_n420_), .C2(new_n422_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n499_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n475_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT98), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n501_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n500_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G78gat), .B(G106gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(G155gat), .A2(G162gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G155gat), .A2(G162gat), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT1), .ZN(new_n521_));
  OR2_X1    g320(.A1(G141gat), .A2(G148gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G141gat), .A2(G148gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT87), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(G155gat), .A2(G162gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT1), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G155gat), .A2(G162gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n524_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(G141gat), .A2(G148gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n530_), .A2(new_n533_), .A3(new_n534_), .A4(new_n523_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n519_), .A2(new_n520_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT3), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT2), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n524_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n526_), .A2(new_n535_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(G228gat), .B(G233gat), .C1(new_n480_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G22gat), .B(G50gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n546_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G228gat), .A2(G233gat), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n435_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n518_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n547_), .A2(new_n553_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n554_), .A3(new_n517_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n514_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G227gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(G71gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n218_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n470_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G127gat), .B(G134gat), .Z(new_n570_));
  XOR2_X1   g369(.A(G113gat), .B(G120gat), .Z(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n569_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G43gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT86), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT30), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT31), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G1gat), .B(G29gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G85gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT0), .B(G57gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G225gat), .A2(G233gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT95), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n526_), .A2(new_n535_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n543_), .A2(new_n536_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT93), .A3(new_n572_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n570_), .B(new_n571_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n544_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n593_), .B2(new_n572_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n544_), .A2(KEYINPUT94), .A3(new_n596_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT4), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT4), .B1(new_n593_), .B2(new_n572_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n590_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n598_), .A2(new_n588_), .A3(new_n601_), .A4(new_n602_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n544_), .A2(KEYINPUT94), .A3(new_n596_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT94), .B1(new_n544_), .B2(new_n596_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n613_), .A2(KEYINPUT96), .A3(new_n588_), .A4(new_n598_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n587_), .B1(new_n607_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT4), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n613_), .B2(new_n598_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n589_), .B1(new_n618_), .B2(new_n605_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(new_n586_), .A3(new_n610_), .A4(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n582_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n564_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT33), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n615_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n626_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n628_), .A2(new_n586_), .A3(new_n619_), .A4(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n502_), .A2(new_n503_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n588_), .B1(new_n618_), .B2(new_n605_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n613_), .A2(new_n598_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n632_), .B(new_n587_), .C1(new_n590_), .C2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n627_), .A2(new_n630_), .A3(new_n631_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n468_), .A2(KEYINPUT32), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n483_), .B2(new_n497_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n506_), .A2(new_n509_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n621_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n563_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n562_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n514_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n582_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n624_), .B1(new_n645_), .B2(KEYINPUT99), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n641_), .A2(new_n563_), .B1(new_n514_), .B2(new_n643_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(new_n582_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n395_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n374_), .A2(new_n375_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n300_), .A3(new_n621_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n291_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n371_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n395_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n322_), .A4(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n660_), .B2(new_n622_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n654_), .A2(new_n655_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n661_), .A3(new_n662_), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n498_), .A2(new_n499_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(KEYINPUT27), .A3(new_n475_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n512_), .B1(new_n511_), .B2(new_n501_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n510_), .C2(new_n475_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n653_), .A2(new_n301_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G8gat), .B1(new_n660_), .B2(new_n514_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT39), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n669_), .A2(KEYINPUT40), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n660_), .B2(new_n581_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT41), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n651_), .A2(G15gat), .A3(new_n581_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1326gat));
  OAI21_X1  g479(.A(G22gat), .B1(new_n660_), .B2(new_n563_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n563_), .A2(G22gat), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT101), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n651_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT102), .ZN(G1327gat));
  INV_X1    g485(.A(new_n291_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n371_), .A2(new_n687_), .A3(new_n322_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n650_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n621_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  INV_X1    g490(.A(new_n322_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n658_), .A2(new_n692_), .A3(new_n659_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT103), .Z(new_n694_));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n564_), .A2(new_n623_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n622_), .A2(new_n562_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n668_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n562_), .B1(new_n635_), .B2(new_n640_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT99), .B(new_n581_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n649_), .A2(new_n697_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n292_), .A2(new_n324_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n695_), .B(new_n696_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n697_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n642_), .A2(new_n644_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n706_), .B2(new_n581_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT43), .B1(new_n708_), .B2(KEYINPUT104), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n704_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n691_), .B1(new_n694_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n693_), .B(KEYINPUT103), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(KEYINPUT44), .C1(new_n704_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n621_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n690_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(new_n689_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(G36gat), .A3(new_n514_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT45), .Z(new_n720_));
  OAI21_X1  g519(.A(G36gat), .B1(new_n714_), .B2(new_n514_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n721_), .A3(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  AOI21_X1  g525(.A(G43gat), .B1(new_n689_), .B2(new_n582_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT105), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n582_), .A2(G43gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n714_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n689_), .B2(new_n562_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n562_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n715_), .B2(new_n733_), .ZN(G1331gat));
  AOI21_X1  g533(.A(new_n659_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n658_), .A2(new_n325_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n621_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n658_), .A2(new_n692_), .A3(new_n659_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n657_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n621_), .B2(KEYINPUT106), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(KEYINPUT106), .B2(new_n743_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n739_), .B1(new_n742_), .B2(new_n745_), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n741_), .B2(new_n514_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT48), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n514_), .A2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n737_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n741_), .B2(new_n581_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n738_), .A2(new_n566_), .A3(new_n582_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n741_), .B2(new_n563_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n563_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n737_), .B2(new_n757_), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n658_), .A2(new_n322_), .A3(new_n659_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n292_), .A2(new_n324_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n696_), .B1(new_n762_), .B2(new_n695_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n708_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n622_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n658_), .A2(new_n322_), .A3(new_n687_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n735_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n203_), .A3(new_n621_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(new_n771_), .ZN(G1336gat));
  OAI21_X1  g571(.A(G92gat), .B1(new_n766_), .B2(new_n514_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n204_), .A3(new_n668_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1337gat));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n218_), .B1(new_n765_), .B2(new_n582_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n234_), .A2(new_n237_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n769_), .A2(new_n778_), .A3(new_n581_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n776_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n777_), .A2(new_n783_), .A3(new_n779_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n786_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(new_n776_), .A3(KEYINPUT51), .A4(new_n784_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1338gat));
  OAI211_X1 g589(.A(new_n562_), .B(new_n759_), .C1(new_n704_), .C2(new_n709_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792_));
  OAI21_X1  g591(.A(G106gat), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT109), .B1(new_n765_), .B2(new_n562_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT52), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n792_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n765_), .A2(KEYINPUT109), .A3(new_n562_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .A4(G106gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n770_), .A2(new_n219_), .A3(new_n562_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n804_), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  NAND2_X1  g605(.A1(new_n582_), .A2(new_n621_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n564_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n388_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT112), .Z(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n380_), .B1(new_n384_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n812_), .B2(new_n384_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n390_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n395_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n336_), .A2(new_n341_), .A3(KEYINPUT55), .A4(new_n342_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT110), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n260_), .A2(new_n261_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n331_), .A2(new_n340_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n340_), .A2(new_n339_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT55), .A4(new_n336_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n342_), .B1(new_n347_), .B2(KEYINPUT12), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n332_), .A2(new_n335_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n341_), .A2(new_n342_), .A3(new_n332_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n334_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n820_), .A2(new_n825_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n352_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n352_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n817_), .B(new_n818_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n816_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n352_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n352_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n818_), .B1(new_n841_), .B2(new_n817_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n687_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n809_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n687_), .C1(new_n836_), .C2(new_n842_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n335_), .B1(new_n347_), .B2(KEYINPUT70), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n339_), .A2(new_n345_), .A3(new_n332_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n823_), .A2(new_n336_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n356_), .B1(new_n850_), .B2(new_n353_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n357_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n815_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT115), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n358_), .A2(new_n855_), .A3(new_n815_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n833_), .A2(new_n834_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n847_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n841_), .A2(KEYINPUT58), .A3(new_n856_), .A4(new_n854_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n703_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n846_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n845_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n817_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT111), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n816_), .A3(new_n835_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866_), .B2(new_n687_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n809_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n322_), .B1(new_n863_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n372_), .B2(new_n395_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n325_), .A2(new_n371_), .A3(KEYINPUT54), .A4(new_n659_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n808_), .B1(new_n869_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G113gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n659_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n692_), .B1(new_n862_), .B2(new_n867_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT116), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n871_), .A2(new_n872_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n692_), .C1(new_n862_), .C2(new_n867_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n880_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n808_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(KEYINPUT59), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n874_), .A2(KEYINPUT59), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n886_), .A2(new_n659_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n877_), .B1(new_n887_), .B2(new_n876_), .ZN(G1340gat));
  NOR2_X1   g687(.A1(new_n658_), .A2(KEYINPUT60), .ZN(new_n889_));
  MUX2_X1   g688(.A(new_n889_), .B(KEYINPUT60), .S(G120gat), .Z(new_n890_));
  NAND2_X1  g689(.A1(new_n875_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n843_), .A2(new_n844_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT114), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n893_), .A2(new_n868_), .A3(new_n846_), .A4(new_n861_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n873_), .B1(new_n894_), .B2(new_n692_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT59), .B1(new_n895_), .B2(new_n884_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n883_), .A2(new_n885_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n371_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT117), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G120gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(KEYINPUT117), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n891_), .B1(new_n900_), .B2(new_n901_), .ZN(G1341gat));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n886_), .B2(new_n322_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n874_), .A2(G127gat), .A3(new_n692_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT118), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n896_), .A2(new_n897_), .A3(new_n322_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G127gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909_));
  INV_X1    g708(.A(new_n905_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n911_), .ZN(G1342gat));
  AOI21_X1  g711(.A(G134gat), .B1(new_n875_), .B2(new_n291_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT119), .B(G134gat), .Z(new_n914_));
  NOR2_X1   g713(.A1(new_n761_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n886_), .B2(new_n915_), .ZN(G1343gat));
  INV_X1    g715(.A(new_n895_), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n668_), .A2(new_n582_), .A3(new_n563_), .A4(new_n622_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n395_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT120), .B(G141gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1344gat));
  NOR2_X1   g721(.A1(new_n919_), .A2(new_n658_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(G148gat), .Z(G1345gat));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n919_), .B2(new_n692_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n917_), .A2(KEYINPUT121), .A3(new_n322_), .A4(new_n918_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n919_), .B2(new_n761_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n687_), .A2(G162gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n919_), .B2(new_n933_), .ZN(G1347gat));
  NOR3_X1   g733(.A1(new_n623_), .A2(new_n562_), .A3(new_n514_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n883_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT22), .B(G169gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n659_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT123), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942_));
  OAI21_X1  g741(.A(G169gat), .B1(new_n942_), .B2(KEYINPUT122), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n935_), .A2(new_n659_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n883_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n942_), .A2(KEYINPUT122), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n947_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n943_), .B(new_n946_), .C1(new_n883_), .C2(new_n944_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n941_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT124), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n952_), .B(new_n941_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1348gat));
  AOI21_X1  g753(.A(G176gat), .B1(new_n937_), .B2(new_n371_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n917_), .A2(new_n935_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n371_), .A2(G176gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(G1349gat));
  NOR3_X1   g757(.A1(new_n936_), .A2(new_n692_), .A3(new_n405_), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n917_), .A2(new_n322_), .A3(new_n935_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n960_), .A2(KEYINPUT125), .ZN(new_n961_));
  AOI21_X1  g760(.A(G183gat), .B1(new_n960_), .B2(KEYINPUT125), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n961_), .B2(new_n962_), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n937_), .A2(new_n291_), .A3(new_n406_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n937_), .A2(new_n703_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(G190gat), .ZN(new_n967_));
  AOI211_X1 g766(.A(KEYINPUT126), .B(new_n445_), .C1(new_n937_), .C2(new_n703_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n964_), .B1(new_n967_), .B2(new_n968_), .ZN(G1351gat));
  NAND3_X1  g768(.A1(new_n668_), .A2(new_n581_), .A3(new_n643_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n895_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(new_n659_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n371_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g774(.A1(new_n971_), .A2(new_n322_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  AND2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n976_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n979_), .B1(new_n976_), .B2(new_n977_), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n971_), .B2(new_n703_), .ZN(new_n982_));
  NOR4_X1   g781(.A1(new_n895_), .A2(G218gat), .A3(new_n687_), .A4(new_n970_), .ZN(new_n983_));
  OR3_X1    g782(.A1(new_n982_), .A2(KEYINPUT127), .A3(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(KEYINPUT127), .B1(new_n982_), .B2(new_n983_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(G1355gat));
endmodule


