//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT21), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT90), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n205_), .B2(G197gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n203_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n211_), .A2(new_n206_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT91), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G211gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(G218gat), .ZN(new_n218_));
  INV_X1    g017(.A(G218gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(G211gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT91), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n202_), .A2(new_n213_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n214_), .A2(new_n215_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT91), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n213_), .A2(new_n202_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n209_), .A2(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G233gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G228gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(G228gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241_));
  NAND3_X1  g040(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G141gat), .ZN(new_n247_));
  INV_X1    g046(.A(G148gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n240_), .A2(new_n242_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n245_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n252_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT29), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n234_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT92), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n234_), .A2(new_n266_), .A3(new_n263_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n211_), .A2(new_n206_), .A3(new_n212_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n216_), .A2(new_n221_), .A3(KEYINPUT21), .A4(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n207_), .B(KEYINPUT89), .ZN(new_n273_));
  OAI22_X1  g072(.A1(new_n223_), .A2(new_n224_), .B1(new_n271_), .B2(KEYINPUT21), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n265_), .A2(new_n267_), .B1(new_n233_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT94), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n262_), .A2(KEYINPUT29), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G22gat), .B(G50gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n277_), .A2(new_n279_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n265_), .A2(new_n267_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n276_), .A2(new_n233_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n287_), .A2(new_n279_), .A3(new_n288_), .ZN(new_n289_));
  OAI22_X1  g088(.A1(new_n280_), .A2(new_n285_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n277_), .A2(new_n279_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n279_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n285_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n291_), .A2(KEYINPUT94), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT24), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT23), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT79), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309_));
  INV_X1    g108(.A(new_n301_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT79), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n304_), .A2(new_n306_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n316_));
  INV_X1    g115(.A(G190gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(KEYINPUT26), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT77), .A3(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT76), .A3(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G183gat), .ZN(new_n327_));
  AOI22_X1  g126(.A1(KEYINPUT25), .A2(new_n327_), .B1(new_n317_), .B2(KEYINPUT26), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n321_), .A2(new_n323_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n300_), .A2(KEYINPUT24), .A3(new_n301_), .A4(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n308_), .A2(new_n315_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT22), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n299_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT81), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n337_), .A3(new_n299_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(G169gat), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n334_), .B2(new_n299_), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT81), .B(G176gat), .C1(new_n333_), .C2(KEYINPUT22), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n298_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n306_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n304_), .A2(new_n306_), .A3(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n339_), .B(new_n342_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n332_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n296_), .B1(new_n349_), .B2(new_n275_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT99), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G169gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n299_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n330_), .B(KEYINPUT97), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n353_), .B(new_n354_), .C1(new_n307_), .C2(new_n347_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n312_), .A2(new_n344_), .A3(new_n331_), .A4(new_n345_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n327_), .A2(KEYINPUT25), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n324_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n319_), .A2(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n317_), .A2(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT96), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT96), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n358_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n356_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n227_), .A2(new_n351_), .A3(new_n355_), .A4(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n355_), .B1(new_n356_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT99), .B1(new_n275_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n350_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n332_), .A2(new_n348_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n296_), .B1(new_n375_), .B2(new_n227_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n275_), .A2(new_n368_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n275_), .A2(KEYINPUT98), .A3(new_n368_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n376_), .A2(new_n377_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT18), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n374_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n295_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n376_), .A2(new_n373_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n227_), .A2(new_n355_), .A3(new_n366_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n350_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n377_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n392_), .B(KEYINPUT27), .C1(new_n386_), .C2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n290_), .A2(new_n294_), .A3(new_n391_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G113gat), .B(G120gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G120gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n252_), .A2(new_n261_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT100), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n252_), .B2(new_n261_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n404_), .A2(new_n406_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n262_), .A2(KEYINPUT100), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n400_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417_));
  INV_X1    g216(.A(new_n251_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n244_), .B1(new_n260_), .B2(KEYINPUT1), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n243_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n259_), .A2(new_n260_), .A3(new_n245_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n413_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n409_), .A3(new_n408_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n417_), .B1(new_n423_), .B2(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n411_), .A2(new_n417_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n400_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n416_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G85gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT4), .B1(new_n412_), .B2(new_n415_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n423_), .A2(new_n414_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n433_), .B1(new_n437_), .B2(new_n400_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n428_), .A2(new_n433_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT31), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n349_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n349_), .B(KEYINPUT30), .ZN(new_n446_));
  INV_X1    g245(.A(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n441_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT84), .B(G15gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(G227gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(G43gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  NAND3_X1  g254(.A1(new_n445_), .A2(new_n448_), .A3(new_n441_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n455_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n449_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n407_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n455_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n459_), .A2(new_n449_), .A3(new_n458_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT85), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n413_), .A3(new_n468_), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n399_), .B(new_n440_), .C1(new_n464_), .C2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n416_), .A2(new_n432_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n427_), .B1(new_n437_), .B2(KEYINPUT4), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT33), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n436_), .A2(new_n438_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n434_), .A2(new_n400_), .A3(new_n425_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n437_), .A2(new_n426_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT101), .B1(new_n478_), .B2(new_n433_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n400_), .B1(new_n423_), .B2(new_n414_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT101), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n432_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n477_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n476_), .A2(new_n392_), .A3(new_n388_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT102), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n389_), .A2(new_n390_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n487_), .A2(KEYINPUT102), .A3(new_n483_), .A4(new_n476_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n374_), .A2(new_n382_), .B1(KEYINPUT32), .B2(new_n386_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n439_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n290_), .A2(new_n294_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT103), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n492_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n500_), .B2(new_n488_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT103), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n398_), .A2(new_n391_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n495_), .A3(new_n439_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n499_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n464_), .A2(new_n469_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n470_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT72), .B(G15gat), .ZN(new_n510_));
  INV_X1    g309(.A(G22gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT73), .B(G8gat), .Z(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n517_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G29gat), .B(G36gat), .Z(new_n522_));
  XOR2_X1   g321(.A(G43gat), .B(G50gat), .Z(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT15), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT75), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n521_), .A2(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n520_), .B(new_n524_), .Z(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G113gat), .B(G141gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n530_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n509_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT6), .ZN(new_n546_));
  INV_X1    g345(.A(G85gat), .ZN(new_n547_));
  INV_X1    g346(.A(G92gat), .ZN(new_n548_));
  OR3_X1    g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT9), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(KEYINPUT9), .ZN(new_n552_));
  INV_X1    g351(.A(G106gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT10), .B(G99gat), .Z(new_n554_));
  AOI211_X1 g353(.A(new_n550_), .B(new_n552_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT65), .ZN(new_n556_));
  AOI211_X1 g355(.A(G99gat), .B(G106gat), .C1(new_n556_), .C2(KEYINPUT7), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n556_), .B2(KEYINPUT7), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n546_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT64), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n551_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT67), .B1(new_n562_), .B2(KEYINPUT8), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT66), .B1(new_n559_), .B2(new_n561_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n546_), .A4(new_n558_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n551_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT8), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n563_), .B2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n564_), .A2(KEYINPUT67), .A3(new_n567_), .A4(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(new_n524_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n573_), .B2(new_n525_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT71), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n544_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n543_), .B(KEYINPUT36), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT68), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT11), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G71gat), .B(G78gat), .Z(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n595_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n599_), .A3(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n521_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n604_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(KEYINPUT17), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n592_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n601_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n573_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n571_), .A2(new_n601_), .A3(new_n572_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT12), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n601_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n619_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n571_), .A2(new_n601_), .A3(new_n572_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n619_), .B1(new_n628_), .B2(new_n624_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n632_), .B(new_n633_), .Z(new_n634_));
  NOR3_X1   g433(.A1(new_n627_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT70), .B1(new_n635_), .B2(KEYINPUT69), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n627_), .A2(new_n630_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n634_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n573_), .A2(new_n625_), .A3(new_n620_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n628_), .A2(new_n624_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(KEYINPUT12), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n629_), .B(new_n638_), .C1(new_n642_), .C2(new_n619_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT69), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT70), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n636_), .A2(new_n639_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n639_), .B1(new_n636_), .B2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n617_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n636_), .A2(new_n646_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n634_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n636_), .A2(new_n639_), .A3(new_n646_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT13), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n616_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n540_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n514_), .A3(new_n440_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT104), .Z(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n505_), .B1(new_n501_), .B2(KEYINPUT103), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n494_), .A2(KEYINPUT103), .A3(new_n496_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n508_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n399_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n507_), .A2(new_n663_), .A3(new_n439_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n585_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n588_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n649_), .A2(new_n654_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n539_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n670_), .A2(new_n614_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n514_), .B1(new_n674_), .B2(new_n440_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT105), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n659_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  NAND3_X1  g477(.A1(new_n656_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n503_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G8gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G8gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n656_), .A2(new_n686_), .A3(new_n507_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT106), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n674_), .A2(new_n507_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G15gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT41), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(KEYINPUT41), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(new_n691_), .A3(new_n692_), .ZN(G1326gat));
  NAND3_X1  g492(.A1(new_n656_), .A2(new_n511_), .A3(new_n495_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n674_), .A2(new_n495_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(G22gat), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(new_n671_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n668_), .A2(new_n614_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n540_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n440_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n590_), .A2(new_n591_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n509_), .B2(new_n592_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n710_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n665_), .A2(new_n708_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n671_), .A2(new_n672_), .A3(new_n614_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT109), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n718_), .B(new_n715_), .C1(new_n711_), .C2(new_n713_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n706_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n715_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT44), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n440_), .A2(G29gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n705_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(new_n706_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n712_), .B1(new_n665_), .B2(new_n708_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n592_), .B(new_n710_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n716_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n718_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n714_), .A2(KEYINPUT109), .A3(new_n716_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n504_), .B1(new_n721_), .B2(KEYINPUT44), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT111), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n737_), .A3(G36gat), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n703_), .A2(G36gat), .A3(new_n504_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(KEYINPUT46), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  NOR3_X1   g544(.A1(new_n703_), .A2(G43gat), .A3(new_n508_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n720_), .A2(new_n507_), .A3(new_n722_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G43gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n748_), .B(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n704_), .B2(new_n495_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n495_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n723_), .B2(new_n753_), .ZN(G1331gat));
  INV_X1    g553(.A(new_n616_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT113), .B1(new_n700_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n671_), .A2(new_n757_), .A3(new_n616_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n756_), .A2(new_n758_), .A3(new_n509_), .A4(new_n672_), .ZN(new_n759_));
  INV_X1    g558(.A(G57gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n440_), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n670_), .A2(new_n672_), .A3(new_n671_), .A4(new_n614_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n440_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n763_), .B2(new_n760_), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n504_), .A2(G64gat), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT114), .Z(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n762_), .A2(new_n503_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G64gat), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT48), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT48), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1333gat));
  INV_X1    g571(.A(G71gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n759_), .A2(new_n773_), .A3(new_n507_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n762_), .A2(new_n507_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G71gat), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1334gat));
  INV_X1    g578(.A(G78gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n759_), .A2(new_n780_), .A3(new_n495_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n762_), .A2(new_n495_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G78gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  NOR4_X1   g585(.A1(new_n509_), .A2(new_n671_), .A3(new_n672_), .A4(new_n701_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n547_), .A3(new_n440_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n649_), .A2(new_n654_), .A3(new_n539_), .A4(new_n614_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT115), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n713_), .B2(new_n711_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(new_n440_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n792_), .B2(new_n547_), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n548_), .A3(new_n503_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n791_), .A2(new_n503_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n548_), .ZN(G1337gat));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n507_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n507_), .A2(new_n554_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n797_), .A2(G99gat), .B1(new_n787_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n799_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n553_), .A3(new_n495_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n791_), .A2(new_n495_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G106gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT52), .B(new_n553_), .C1(new_n791_), .C2(new_n495_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  AND4_X1   g609(.A1(new_n810_), .A2(new_n671_), .A3(new_n539_), .A4(new_n755_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n655_), .B2(new_n539_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n623_), .A2(new_n626_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n623_), .A2(new_n816_), .A3(new_n626_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n619_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n819_), .B(new_n820_), .C1(new_n642_), .C2(new_n619_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT55), .B1(new_n627_), .B2(KEYINPUT117), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n634_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT121), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n634_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n823_), .A2(new_n828_), .A3(KEYINPUT56), .A4(new_n634_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n527_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n536_), .B1(new_n531_), .B2(new_n529_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(new_n537_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n635_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n830_), .A2(KEYINPUT58), .A3(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n708_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n827_), .A2(new_n845_), .A3(new_n824_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n539_), .A2(new_n635_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n823_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n634_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n647_), .A2(new_n648_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n837_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n846_), .A2(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n844_), .B1(new_n852_), .B2(new_n668_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n824_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n855_), .A2(new_n826_), .A3(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n847_), .A2(new_n848_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n843_), .A2(new_n853_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n813_), .B1(new_n860_), .B2(new_n614_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n507_), .A2(new_n663_), .A3(new_n440_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT122), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n672_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n852_), .A2(new_n844_), .A3(new_n668_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n858_), .B2(new_n669_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n615_), .B1(new_n870_), .B2(new_n843_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT59), .B(new_n863_), .C1(new_n871_), .C2(new_n813_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n539_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n867_), .B1(new_n875_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n671_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n865_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n671_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n877_), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n872_), .A2(new_n874_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n615_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n865_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n615_), .A2(new_n882_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n614_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n890_));
  OAI221_X1 g689(.A(new_n889_), .B1(new_n885_), .B2(new_n886_), .C1(new_n890_), .C2(new_n882_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(G1342gat));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n865_), .A2(new_n893_), .A3(new_n668_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n592_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1343gat));
  NOR2_X1   g695(.A1(new_n507_), .A2(new_n496_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(new_n503_), .A3(new_n439_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n861_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n861_), .A2(KEYINPUT124), .A3(new_n900_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n672_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g704(.A(new_n700_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g706(.A(new_n615_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  NAND2_X1  g709(.A1(new_n708_), .A2(G162gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT125), .Z(new_n912_));
  INV_X1    g711(.A(new_n903_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n901_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n668_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n915_));
  INV_X1    g714(.A(G162gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1347gat));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n507_), .A2(new_n496_), .A3(new_n503_), .A4(new_n439_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n861_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n539_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n918_), .B1(new_n922_), .B2(new_n298_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n352_), .ZN(new_n924_));
  OAI211_X1 g723(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(new_n539_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  NAND2_X1  g725(.A1(new_n920_), .A2(new_n700_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n921_), .A2(new_n614_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(G183gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n929_), .B2(new_n358_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n921_), .B2(new_n592_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n362_), .A2(new_n364_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n920_), .A2(new_n933_), .A3(new_n668_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(G1351gat));
  INV_X1    g734(.A(new_n861_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n898_), .A2(new_n504_), .A3(new_n440_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n539_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n203_), .ZN(G1352gat));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n671_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(G204gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1353gat));
  INV_X1    g742(.A(new_n938_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n615_), .B1(new_n945_), .B2(new_n217_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT127), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n944_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n945_), .A2(new_n217_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n938_), .B2(new_n592_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n668_), .A2(new_n219_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n938_), .B2(new_n952_), .ZN(G1355gat));
endmodule


