//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(G8gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G8gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT75), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n204_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n207_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G1gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G8gat), .A3(new_n208_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G29gat), .B(G36gat), .Z(new_n215_));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216_));
  XOR2_X1   g015(.A(new_n215_), .B(new_n216_), .Z(new_n217_));
  AND3_X1   g016(.A1(new_n211_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n219_));
  OAI211_X1 g018(.A(G229gat), .B(G233gat), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G141gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT78), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n211_), .A2(new_n214_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n217_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n217_), .B(KEYINPUT15), .Z(new_n231_));
  NAND3_X1  g030(.A1(new_n211_), .A2(new_n214_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT77), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n220_), .A2(new_n227_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n227_), .B1(new_n220_), .B2(new_n236_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT79), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G78gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(G57gat), .B(G64gat), .Z(new_n245_));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n246_), .B2(new_n245_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n244_), .A3(KEYINPUT11), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT10), .B(G99gat), .Z(new_n256_));
  INV_X1    g055(.A(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G85gat), .B(G92gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT9), .ZN(new_n260_));
  INV_X1    g059(.A(G85gat), .ZN(new_n261_));
  INV_X1    g060(.A(G92gat), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT9), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G99gat), .A2(G106gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT6), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n258_), .A2(new_n260_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT8), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n270_));
  NOR2_X1   g069(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n270_), .A2(new_n271_), .B1(G99gat), .B2(G106gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n265_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT65), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT65), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n269_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n273_), .B1(new_n283_), .B2(new_n274_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n273_), .A2(new_n274_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n280_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n272_), .A2(KEYINPUT66), .A3(new_n275_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n265_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n259_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n268_), .B1(new_n289_), .B2(KEYINPUT67), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n291_), .A3(new_n259_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n279_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n254_), .B(new_n255_), .C1(new_n267_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(KEYINPUT67), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(KEYINPUT8), .A3(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n279_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n267_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n251_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT12), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT69), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n253_), .B1(new_n298_), .B2(new_n251_), .ZN(new_n303_));
  AND2_X1   g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n298_), .B2(new_n251_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n294_), .A2(new_n302_), .A3(new_n303_), .A4(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n298_), .A2(new_n251_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n251_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n293_), .A2(new_n308_), .A3(new_n267_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n304_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G120gat), .B(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT5), .B(G176gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  AND3_X1   g114(.A1(new_n306_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT13), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT13), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G64gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(new_n262_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n312_), .A2(G197gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n223_), .A2(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G218gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G211gat), .ZN(new_n332_));
  INV_X1    g131(.A(G211gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G218gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n332_), .A2(new_n334_), .A3(KEYINPUT90), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT90), .B1(new_n332_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n330_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n312_), .B2(G197gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n223_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n327_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n337_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n329_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n333_), .A2(G218gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n331_), .A2(G211gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n332_), .A2(new_n334_), .A3(KEYINPUT90), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n350_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(KEYINPUT91), .A3(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n348_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n357_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(new_n359_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n347_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n367_), .A2(KEYINPUT24), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT80), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT23), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n367_), .A2(KEYINPUT24), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT25), .B(G183gat), .Z(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT26), .B(G190gat), .Z(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n370_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(G176gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G169gat), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n372_), .A2(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n368_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n361_), .A2(new_n359_), .A3(new_n349_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT92), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n346_), .B1(new_n388_), .B2(new_n362_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT93), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n366_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n364_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(KEYINPUT94), .ZN(new_n394_));
  AOI211_X1 g193(.A(new_n369_), .B(new_n378_), .C1(new_n375_), .C2(KEYINPUT97), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n375_), .A2(KEYINPUT97), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n368_), .B(KEYINPUT98), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n395_), .A2(new_n396_), .B1(new_n384_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n399_), .A3(KEYINPUT20), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n380_), .A2(new_n385_), .ZN(new_n404_));
  AOI211_X1 g203(.A(new_n365_), .B(new_n346_), .C1(new_n388_), .C2(new_n362_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n388_), .A2(new_n362_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT93), .B1(new_n406_), .B2(new_n347_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n395_), .A2(new_n396_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n384_), .A2(new_n397_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n413_), .B2(new_n364_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n326_), .B1(new_n403_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n402_), .B1(new_n398_), .B2(new_n389_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n391_), .A2(KEYINPUT20), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n409_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n416_), .B1(new_n326_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(KEYINPUT1), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT84), .B(new_n423_), .C1(new_n424_), .C2(KEYINPUT1), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n427_), .B(new_n428_), .C1(KEYINPUT1), .C2(new_n423_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G141gat), .B(G148gat), .Z(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n423_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n432_), .A2(new_n424_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n432_), .B2(new_n424_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT3), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(G141gat), .B2(G148gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n436_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT87), .B(new_n436_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n431_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G127gat), .B(G134gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G120gat), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n455_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n453_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n456_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n459_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI211_X1 g263(.A(new_n464_), .B(new_n431_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT4), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n431_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n442_), .A2(new_n445_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT85), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT87), .B1(new_n473_), .B2(new_n436_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n452_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n460_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT4), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n466_), .A2(new_n468_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT0), .ZN(new_n483_));
  INV_X1    g282(.A(G57gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n261_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n478_), .B1(new_n476_), .B2(new_n464_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n467_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT99), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n481_), .A2(KEYINPUT99), .A3(new_n488_), .A4(new_n486_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n481_), .A2(new_n488_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n491_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n422_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n386_), .B1(new_n366_), .B2(new_n390_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT20), .B1(new_n398_), .B2(new_n389_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n402_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n325_), .A3(new_n418_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n486_), .B1(new_n487_), .B2(new_n467_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n466_), .A2(new_n480_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n467_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n325_), .B1(new_n500_), .B2(new_n418_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n502_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT33), .B1(new_n493_), .B2(new_n494_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509_));
  AOI211_X1 g308(.A(new_n509_), .B(new_n486_), .C1(new_n481_), .C2(new_n488_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n497_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n476_), .A2(KEYINPUT29), .ZN(new_n514_));
  XOR2_X1   g313(.A(G22gat), .B(G50gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT28), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n514_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G78gat), .B(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n476_), .A2(KEYINPUT29), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n366_), .A3(new_n522_), .A4(new_n390_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n393_), .A2(new_n394_), .B1(KEYINPUT29), .B2(new_n476_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n520_), .B(new_n523_), .C1(new_n524_), .C2(new_n522_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n389_), .A2(KEYINPUT94), .ZN(new_n526_));
  AOI211_X1 g325(.A(new_n392_), .B(new_n346_), .C1(new_n388_), .C2(new_n362_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n521_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n522_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n520_), .B1(new_n530_), .B2(new_n523_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n525_), .B1(new_n531_), .B2(KEYINPUT95), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n530_), .A2(new_n533_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n518_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n525_), .A2(KEYINPUT96), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n523_), .B1(new_n524_), .B2(new_n522_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n519_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n530_), .A2(new_n539_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(new_n518_), .A3(new_n538_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G99gat), .Z(new_n543_));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G15gat), .B(G43gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n404_), .A2(KEYINPUT30), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n386_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT81), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n477_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n477_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n550_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n535_), .A2(new_n542_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n513_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n525_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n534_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n517_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n561_), .A2(new_n563_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n541_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n564_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n501_), .A2(KEYINPUT27), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n325_), .B(KEYINPUT100), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n403_), .B2(new_n415_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n578_));
  INV_X1    g377(.A(new_n325_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n580_), .B2(new_n501_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n577_), .A2(new_n496_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n573_), .A3(new_n582_), .ZN(new_n583_));
  AOI211_X1 g382(.A(new_n243_), .B(new_n321_), .C1(new_n566_), .C2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n231_), .B1(new_n293_), .B2(new_n267_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n288_), .A2(new_n291_), .A3(new_n259_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n291_), .B1(new_n288_), .B2(new_n259_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n268_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n266_), .B(new_n229_), .C1(new_n588_), .C2(new_n279_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT35), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT70), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n595_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(KEYINPUT35), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n592_), .B1(new_n298_), .B2(new_n229_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(new_n585_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT71), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT72), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n601_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(KEYINPUT73), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n607_), .B(new_n612_), .C1(KEYINPUT73), .C2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n228_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n300_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n252_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n625_));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G183gat), .B(G211gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n623_), .A2(KEYINPUT17), .A3(new_n624_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n622_), .A2(new_n251_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n621_), .A2(new_n308_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n629_), .B(KEYINPUT17), .Z(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n619_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n584_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n204_), .A3(new_n496_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n566_), .A2(new_n583_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n613_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n239_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n644_), .A2(new_n321_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n204_), .B1(new_n646_), .B2(new_n496_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n640_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n639_), .B2(new_n638_), .ZN(G1324gat));
  INV_X1    g448(.A(new_n577_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n581_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n202_), .B1(new_n646_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT39), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n637_), .A2(new_n203_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n646_), .B2(new_n564_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n637_), .A2(new_n658_), .A3(new_n564_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n535_), .A2(new_n542_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n646_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT102), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n637_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n635_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n613_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n584_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n496_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n615_), .A2(new_n676_), .A3(new_n617_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n566_), .B2(new_n583_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n572_), .A2(new_n573_), .A3(new_n582_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n496_), .A2(new_n422_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n572_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n615_), .A2(KEYINPUT103), .A3(new_n617_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT103), .B1(new_n615_), .B2(new_n617_), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n679_), .A2(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n678_), .B1(new_n684_), .B2(KEYINPUT43), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n321_), .A2(new_n671_), .A3(new_n645_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n675_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT104), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n618_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n615_), .A2(KEYINPUT103), .A3(new_n617_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n676_), .B1(new_n693_), .B2(new_n641_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n686_), .B1(new_n694_), .B2(new_n678_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n675_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n689_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n686_), .C1(new_n694_), .C2(new_n678_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(G29gat), .A3(new_n496_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n674_), .B1(new_n698_), .B2(new_n700_), .ZN(G1328gat));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n652_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n650_), .A2(KEYINPUT106), .A3(new_n651_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n673_), .A2(new_n702_), .A3(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n699_), .A2(new_n652_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n689_), .B2(new_n697_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G36gat), .B1(new_n711_), .B2(KEYINPUT105), .ZN(new_n712_));
  INV_X1    g511(.A(new_n710_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n688_), .A2(KEYINPUT104), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n696_), .B1(new_n695_), .B2(new_n675_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT105), .B(new_n713_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n709_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT46), .B(new_n709_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NAND4_X1  g521(.A1(new_n698_), .A2(G43gat), .A3(new_n564_), .A4(new_n699_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n673_), .A2(new_n564_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(G43gat), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n673_), .B2(new_n665_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n699_), .A2(G50gat), .A3(new_n665_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n698_), .B2(new_n728_), .ZN(G1331gat));
  INV_X1    g528(.A(new_n496_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n641_), .A2(new_n645_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT107), .ZN(new_n733_));
  INV_X1    g532(.A(new_n321_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n636_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n730_), .B1(new_n736_), .B2(KEYINPUT108), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(KEYINPUT108), .B2(new_n736_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n243_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n644_), .A2(new_n734_), .A3(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n730_), .A2(new_n484_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n738_), .A2(new_n484_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n740_), .B2(new_n707_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT110), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n744_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n707_), .A2(new_n743_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n736_), .B2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n740_), .B2(new_n564_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT49), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n564_), .A2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n736_), .B2(new_n753_), .ZN(G1334gat));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n740_), .B2(new_n665_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT50), .Z(new_n757_));
  NAND2_X1  g556(.A1(new_n665_), .A2(new_n755_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n736_), .B2(new_n758_), .ZN(G1335gat));
  NOR3_X1   g558(.A1(new_n734_), .A2(new_n671_), .A3(new_n239_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n694_), .B2(new_n678_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n762_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n730_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n735_), .A2(new_n672_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n261_), .A3(new_n496_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n706_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n262_), .A3(new_n652_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1337gat));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n256_), .A3(new_n564_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n571_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n774_));
  INV_X1    g573(.A(G99gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n257_), .A3(new_n665_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G106gat), .B1(new_n761_), .B2(new_n664_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT52), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT52), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g582(.A1(new_n652_), .A2(new_n571_), .A3(new_n730_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n316_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n302_), .A2(new_n303_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n294_), .A4(new_n305_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n298_), .A2(new_n251_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n294_), .A2(new_n302_), .A3(new_n303_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n304_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n306_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n315_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n315_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n791_), .A2(new_n306_), .B1(new_n789_), .B2(new_n304_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n787_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n785_), .B1(new_n795_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n225_), .B1(new_n220_), .B2(new_n236_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n235_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n230_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n224_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n318_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n642_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n793_), .A2(new_n797_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n315_), .B1(new_n799_), .B2(new_n787_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(KEYINPUT56), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n813_), .B2(new_n785_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n642_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n810_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n793_), .A2(new_n794_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n796_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n811_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n800_), .A2(KEYINPUT112), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n806_), .A2(new_n316_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n824_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n619_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n671_), .B1(new_n817_), .B2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n739_), .A2(new_n321_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n636_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n636_), .B2(new_n831_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n664_), .B(new_n784_), .C1(new_n830_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT113), .ZN(new_n837_));
  INV_X1    g636(.A(new_n835_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n824_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n823_), .B2(new_n824_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n618_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n815_), .B1(new_n814_), .B2(new_n642_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n635_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n838_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n664_), .A4(new_n784_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n837_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G113gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n239_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n846_), .A2(new_n853_), .A3(new_n664_), .A4(new_n784_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n243_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n851_), .A2(new_n856_), .ZN(G1340gat));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n734_), .B2(G120gat), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n837_), .A2(new_n848_), .A3(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n852_), .A2(new_n854_), .A3(new_n321_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G120gat), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n855_), .A2(new_n865_), .A3(new_n635_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n837_), .A2(new_n848_), .A3(new_n671_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n865_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT114), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n870_), .A3(new_n865_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n866_), .B1(new_n869_), .B2(new_n871_), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n849_), .A2(new_n642_), .ZN(new_n873_));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n855_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n619_), .A2(G134gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT115), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n873_), .A2(new_n874_), .B1(new_n875_), .B2(new_n877_), .ZN(G1343gat));
  NAND3_X1  g677(.A1(new_n704_), .A2(new_n496_), .A3(new_n705_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n664_), .A2(new_n564_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n879_), .A2(new_n881_), .A3(KEYINPUT116), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT116), .B1(new_n879_), .B2(new_n881_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n838_), .B2(new_n845_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n239_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT117), .B(G141gat), .Z(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n321_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT118), .B(G148gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1345gat));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n885_), .A2(new_n894_), .A3(new_n671_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n884_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n671_), .C1(new_n830_), .C2(new_n835_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT119), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n893_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n895_), .A2(new_n898_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT120), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n892_), .A3(new_n900_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n885_), .A2(new_n642_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n909_), .A2(KEYINPUT121), .A3(G162gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n909_), .B2(G162gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n693_), .A2(G162gat), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n885_), .B2(new_n912_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n830_), .A2(new_n835_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n665_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n706_), .A2(new_n571_), .A3(new_n496_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917_), .B2(new_n645_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  OAI211_X1 g719(.A(KEYINPUT62), .B(G169gat), .C1(new_n917_), .C2(new_n645_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n917_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n383_), .A3(new_n239_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(new_n921_), .A3(new_n923_), .ZN(G1348gat));
  OAI211_X1 g723(.A(new_n922_), .B(new_n321_), .C1(KEYINPUT122), .C2(G176gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT122), .B(G176gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n917_), .B2(new_n734_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1349gat));
  AOI21_X1  g727(.A(G183gat), .B1(new_n922_), .B2(new_n671_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n917_), .A2(new_n635_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n376_), .B2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n917_), .B2(new_n618_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n613_), .A2(new_n377_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n917_), .B2(new_n933_), .ZN(G1351gat));
  NOR3_X1   g733(.A1(new_n706_), .A2(new_n496_), .A3(new_n881_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n914_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n938_), .B(new_n935_), .C1(new_n830_), .C2(new_n835_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n645_), .B1(KEYINPUT124), .B2(new_n223_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n223_), .A2(KEYINPUT124), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT125), .Z(new_n944_));
  XNOR2_X1  g743(.A(new_n942_), .B(new_n944_), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n940_), .A2(new_n321_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g746(.A(KEYINPUT63), .B(G211gat), .Z(new_n948_));
  AOI21_X1  g747(.A(new_n938_), .B1(new_n846_), .B2(new_n935_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n939_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n671_), .B(new_n948_), .C1(new_n949_), .C2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n949_), .A2(new_n950_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n635_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n940_), .A2(KEYINPUT126), .A3(new_n671_), .A4(new_n948_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n953_), .A2(new_n956_), .A3(new_n957_), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n955_), .B2(new_n618_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n940_), .A2(new_n331_), .A3(new_n642_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1355gat));
endmodule


