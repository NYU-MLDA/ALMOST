//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G15gat), .A2(G22gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(G15gat), .A2(G22gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT79), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n208_), .A2(new_n207_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n206_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n203_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(KEYINPUT79), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n211_), .A3(new_n206_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n202_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G29gat), .B(G36gat), .Z(new_n219_));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G29gat), .B(G36gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n225_), .B(KEYINPUT83), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n214_), .A2(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT84), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n225_), .B(new_n237_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n218_), .A2(new_n238_), .A3(KEYINPUT85), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT85), .B1(new_n218_), .B2(new_n238_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n233_), .A3(new_n240_), .A4(new_n228_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n232_), .A2(new_n242_), .A3(new_n234_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n236_), .A2(new_n241_), .A3(new_n243_), .A4(new_n247_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT86), .B1(new_n249_), .B2(new_n250_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT65), .B(G85gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT9), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(G92gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(G85gat), .A2(G92gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G85gat), .A2(G92gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT9), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT66), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT67), .B(KEYINPUT6), .Z(new_n262_));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G99gat), .A3(G106gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n256_), .A2(new_n268_), .A3(new_n259_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT10), .B(G99gat), .Z(new_n270_));
  INV_X1    g069(.A(G106gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n261_), .A2(new_n267_), .A3(new_n269_), .A4(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G99gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT7), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n274_), .B(new_n271_), .C1(new_n275_), .C2(KEYINPUT68), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(KEYINPUT7), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n275_), .A2(new_n274_), .A3(new_n271_), .A4(KEYINPUT68), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n264_), .A2(new_n266_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT8), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n257_), .A2(new_n258_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n273_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n294_), .A2(KEYINPUT69), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(KEYINPUT69), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n285_), .B(new_n293_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n280_), .A2(new_n282_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT8), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n272_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n268_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n299_), .A2(new_n300_), .B1(new_n269_), .B2(new_n303_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(new_n304_), .A2(new_n292_), .B1(KEYINPUT69), .B2(new_n294_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n273_), .B(new_n292_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT64), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT70), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n297_), .B(new_n305_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n308_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n304_), .A2(new_n292_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n306_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G176gat), .B(G204gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(KEYINPUT71), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n326_), .A2(new_n327_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(KEYINPUT90), .A2(G183gat), .A3(G190gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT90), .B1(G183gat), .B2(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT23), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT87), .B(G183gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n336_), .B(new_n339_), .C1(G190gat), .C2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G169gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n348_), .A2(KEYINPUT24), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT88), .B1(new_n352_), .B2(G190gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G190gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(KEYINPUT88), .ZN(new_n355_));
  NOR2_X1   g154(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n340_), .B2(KEYINPUT25), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n351_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n338_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n348_), .A2(new_n349_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(KEYINPUT24), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n344_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n367_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(G15gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT30), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n371_), .B(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G78gat), .B(G106gat), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT97), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT93), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT2), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n381_), .A2(new_n383_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT91), .B(KEYINPUT3), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT92), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n393_), .B(new_n390_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n386_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(KEYINPUT1), .B2(new_n399_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n399_), .A2(KEYINPUT1), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT94), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n410_));
  AOI211_X1 g209(.A(new_n410_), .B(new_n407_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n415_), .A2(KEYINPUT21), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT21), .B1(new_n415_), .B2(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n414_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(KEYINPUT21), .A3(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(G228gat), .B2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n379_), .B1(new_n413_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n403_), .A2(new_n408_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n410_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n403_), .A2(KEYINPUT94), .A3(new_n408_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT29), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT97), .A3(new_n424_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G228gat), .ZN(new_n433_));
  INV_X1    g232(.A(G233gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(KEYINPUT29), .ZN(new_n435_));
  INV_X1    g234(.A(new_n423_), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n433_), .B(new_n434_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n378_), .B1(new_n432_), .B2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n377_), .B(new_n437_), .C1(new_n426_), .C2(new_n431_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G22gat), .B(G50gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT96), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n428_), .A2(new_n429_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n412_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n412_), .B(new_n444_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n409_), .A2(new_n411_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n443_), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n451_));
  INV_X1    g250(.A(new_n441_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n439_), .A2(new_n440_), .A3(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n446_), .A2(new_n448_), .A3(new_n441_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n451_), .B2(new_n447_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n413_), .A2(new_n379_), .A3(new_n425_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT97), .B1(new_n430_), .B2(new_n424_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n438_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n377_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n432_), .A2(new_n378_), .A3(new_n438_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n458_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n455_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT18), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n423_), .B(new_n344_), .C1(new_n358_), .C2(new_n363_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT20), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n361_), .B2(new_n475_), .ZN(new_n476_));
  AOI211_X1 g275(.A(KEYINPUT101), .B(new_n474_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n343_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n339_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n337_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT90), .A2(G183gat), .A3(G190gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n479_), .B1(new_n483_), .B2(KEYINPUT23), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n348_), .A2(new_n349_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n348_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT25), .B(G183gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n354_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT100), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n485_), .A2(new_n486_), .B1(new_n354_), .B2(new_n490_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT100), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n489_), .A4(new_n484_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n478_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n472_), .B1(new_n436_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT19), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT98), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT102), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(new_n496_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n343_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n361_), .A2(new_n475_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT101), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n361_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n436_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n471_), .A2(KEYINPUT20), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT102), .ZN(new_n512_));
  INV_X1    g311(.A(new_n501_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n502_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n478_), .A2(new_n423_), .A3(new_n493_), .A4(new_n496_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n364_), .B2(new_n436_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n500_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n470_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n469_), .B(new_n522_), .C1(new_n502_), .C2(new_n514_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G29gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G85gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT0), .B(G57gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT4), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n428_), .A2(new_n429_), .A3(new_n370_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n427_), .A2(new_n370_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT4), .B1(new_n450_), .B2(new_n370_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n533_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n536_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n529_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT103), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n536_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n531_), .A2(new_n533_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n528_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n531_), .A2(new_n530_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n532_), .B1(new_n450_), .B2(new_n370_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n530_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n536_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n545_), .B(new_n548_), .C1(new_n549_), .C2(new_n530_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n528_), .B1(new_n552_), .B2(new_n539_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n553_), .B2(KEYINPUT33), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT103), .B1(new_n553_), .B2(KEYINPUT33), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n524_), .A2(new_n544_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n478_), .A2(new_n423_), .A3(new_n492_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n518_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n500_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n515_), .A2(new_n520_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n537_), .A2(new_n540_), .A3(new_n529_), .ZN(new_n564_));
  OAI221_X1 g363(.A(new_n562_), .B1(new_n563_), .B2(new_n561_), .C1(new_n564_), .C2(new_n553_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n465_), .B1(new_n556_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT27), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n560_), .A2(new_n469_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT27), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT104), .B1(new_n523_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n515_), .A2(new_n470_), .A3(new_n520_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT104), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT27), .A4(new_n569_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n564_), .A2(new_n553_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n454_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n462_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n376_), .B1(new_n566_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n575_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n465_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n376_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n576_), .A4(new_n584_), .ZN(new_n585_));
  AOI211_X1 g384(.A(new_n253_), .B(new_n333_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n238_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n285_), .A2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n273_), .B(new_n225_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT35), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT75), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(KEYINPUT35), .B2(new_n592_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n593_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n589_), .A2(new_n590_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT76), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n589_), .A2(new_n601_), .A3(new_n590_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT73), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT74), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n607_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n589_), .A2(new_n590_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n594_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n603_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n587_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n609_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT77), .B1(new_n612_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT77), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n611_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n600_), .A2(new_n602_), .B1(new_n613_), .B2(new_n594_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n615_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n617_), .A2(new_n625_), .ZN(new_n626_));
  OAI221_X1 g425(.A(new_n615_), .B1(new_n616_), .B2(new_n587_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n292_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n230_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G127gat), .B(G155gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n636_));
  NOR3_X1   g435(.A1(new_n631_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n635_), .B(KEYINPUT17), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT81), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(KEYINPUT81), .A3(new_n638_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n637_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n628_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT82), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n586_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT105), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n576_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n204_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n625_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n643_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n586_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n576_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n655_), .A3(new_n660_), .ZN(G1324gat));
  OAI21_X1  g460(.A(G8gat), .B1(new_n659_), .B2(new_n582_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n575_), .A2(new_n205_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n649_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n665_), .B(new_n666_), .Z(G1325gat));
  NOR3_X1   g466(.A1(new_n649_), .A2(G15gat), .A3(new_n376_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT107), .Z(new_n669_));
  OAI21_X1  g468(.A(G15gat), .B1(new_n659_), .B2(new_n376_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT41), .Z(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1326gat));
  OAI21_X1  g471(.A(G22gat), .B1(new_n659_), .B2(new_n583_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n583_), .A2(G22gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT108), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n649_), .B2(new_n676_), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n625_), .A2(new_n643_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n586_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G29gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n651_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n333_), .A2(new_n253_), .A3(new_n643_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n626_), .A2(KEYINPUT109), .A3(new_n627_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n581_), .A2(new_n585_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n628_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n628_), .B(new_n684_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n682_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n651_), .A3(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT110), .B1(new_n694_), .B2(G29gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n681_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n575_), .A3(new_n693_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT111), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n692_), .A2(new_n700_), .A3(new_n575_), .A4(new_n693_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n699_), .A2(G36gat), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n679_), .A2(new_n703_), .A3(new_n575_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NAND2_X1  g504(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n702_), .A2(new_n705_), .B1(KEYINPUT112), .B2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n698_), .A2(KEYINPUT111), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n701_), .A2(G36gat), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT112), .B(new_n705_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT113), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1329gat));
  NAND2_X1  g512(.A1(new_n692_), .A2(new_n693_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G43gat), .B1(new_n714_), .B2(new_n376_), .ZN(new_n715_));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n679_), .A2(new_n716_), .A3(new_n584_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n714_), .B2(new_n583_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n583_), .A2(G50gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT114), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n679_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1331gat));
  NOR2_X1   g523(.A1(KEYINPUT116), .A2(G57gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n253_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n726_), .B(new_n332_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n658_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n576_), .A2(KEYINPUT116), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n725_), .B(new_n728_), .C1(G57gat), .C2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n645_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT115), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(KEYINPUT115), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n651_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n730_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n728_), .B2(new_n582_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n582_), .A2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n731_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n728_), .B2(new_n376_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n376_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n731_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n728_), .B2(new_n583_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n583_), .A2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n731_), .B2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n727_), .A2(new_n678_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n651_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n688_), .A2(new_n689_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n726_), .A2(new_n332_), .A3(new_n643_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n651_), .A2(new_n254_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  INV_X1    g556(.A(G92gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(new_n758_), .A3(new_n575_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n575_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n761_), .B2(new_n758_), .ZN(G1337gat));
  AND3_X1   g561(.A1(new_n751_), .A2(new_n270_), .A3(new_n584_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n755_), .A2(new_n584_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G99gat), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT51), .Z(G1338gat));
  OAI211_X1 g565(.A(new_n465_), .B(new_n754_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G106gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT52), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n751_), .A2(new_n271_), .A3(new_n465_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1339gat));
  NOR3_X1   g572(.A1(new_n657_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n332_), .A3(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n628_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT118), .B1(new_n774_), .B2(new_n332_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT119), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n332_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n628_), .A4(new_n775_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(KEYINPUT54), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT119), .B(new_n785_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n313_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n249_), .A2(new_n250_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT86), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n250_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n305_), .A2(new_n297_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n314_), .B1(new_n794_), .B2(new_n316_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n313_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n305_), .A2(new_n297_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(KEYINPUT55), .C1(new_n312_), .C2(new_n310_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT120), .B(new_n314_), .C1(new_n794_), .C2(new_n316_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n797_), .A2(new_n799_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n321_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n321_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n793_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n247_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT121), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n239_), .A2(new_n240_), .A3(new_n228_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n233_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n250_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n656_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n250_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n788_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT122), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n628_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n805_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n321_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(KEYINPUT58), .A4(new_n815_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n819_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n812_), .A2(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n813_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n657_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n376_), .B1(new_n787_), .B2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n575_), .A2(new_n465_), .A3(new_n576_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n726_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n830_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n253_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n838_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n332_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n831_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n332_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n831_), .A2(new_n845_), .A3(new_n643_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n657_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n835_), .B2(new_n625_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(KEYINPUT123), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n687_), .A2(G134gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n850_), .A2(KEYINPUT123), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .ZN(G1343gat));
  AOI21_X1  g654(.A(new_n584_), .B1(new_n787_), .B2(new_n828_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(new_n465_), .A3(new_n651_), .A4(new_n582_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n253_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n332_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g660(.A1(new_n857_), .A2(new_n657_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n857_), .B2(new_n628_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n625_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n857_), .B2(new_n866_), .ZN(G1347gat));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n582_), .A2(new_n651_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n465_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n812_), .A2(KEYINPUT57), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n873_), .B(new_n656_), .C1(new_n806_), .C2(new_n811_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n643_), .B1(new_n875_), .B2(new_n825_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n784_), .A2(new_n786_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n584_), .B(new_n871_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n726_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n868_), .B1(new_n880_), .B2(G169gat), .ZN(new_n881_));
  AOI211_X1 g680(.A(KEYINPUT62), .B(new_n346_), .C1(new_n879_), .C2(new_n726_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n829_), .B2(new_n871_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n878_), .A2(KEYINPUT124), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT22), .B(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n726_), .A2(new_n887_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n881_), .A2(new_n882_), .B1(new_n886_), .B2(new_n888_), .ZN(G1348gat));
  OAI21_X1  g688(.A(G176gat), .B1(new_n878_), .B2(new_n332_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n333_), .A2(new_n347_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n886_), .B2(new_n891_), .ZN(G1349gat));
  OR2_X1    g691(.A1(new_n657_), .A2(new_n490_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n878_), .A2(KEYINPUT124), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n787_), .A2(new_n828_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n895_), .A2(new_n883_), .A3(new_n584_), .A4(new_n871_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n878_), .A2(new_n657_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n340_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  OR3_X1    g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g702(.A(new_n687_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT126), .B1(new_n904_), .B2(G190gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n628_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  INV_X1    g706(.A(G190gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n656_), .A2(new_n354_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n905_), .A2(new_n909_), .B1(new_n886_), .B2(new_n910_), .ZN(G1351gat));
  NOR2_X1   g710(.A1(new_n870_), .A2(new_n583_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n856_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n253_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT127), .B(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n332_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g717(.A1(new_n913_), .A2(new_n657_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n919_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT63), .B(G211gat), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(G1354gat));
  OAI21_X1  g721(.A(G218gat), .B1(new_n913_), .B2(new_n628_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n625_), .A2(G218gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n913_), .B2(new_n924_), .ZN(G1355gat));
endmodule


