//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  INV_X1    g006(.A(G43gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(G50gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT76), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(KEYINPUT14), .C1(new_n211_), .C2(new_n212_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G1gat), .B(G8gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n219_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n210_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT81), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G50gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n209_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT15), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n210_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n223_), .B(new_n226_), .C1(new_n232_), .C2(new_n222_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n210_), .A2(new_n222_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n224_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n206_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n206_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n222_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n234_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n239_), .C1(new_n241_), .C2(new_n226_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n242_), .A3(KEYINPUT82), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n244_), .B(new_n206_), .C1(new_n233_), .C2(new_n236_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT10), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(G99gat), .ZN(new_n250_));
  INV_X1    g049(.A(G99gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT10), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n248_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G85gat), .ZN(new_n257_));
  INV_X1    g056(.A(G92gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n254_), .A2(new_n259_), .A3(new_n255_), .A4(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n253_), .A2(new_n256_), .A3(new_n261_), .A4(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT8), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n259_), .A2(new_n255_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n251_), .A2(new_n248_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n266_), .B(new_n267_), .C1(new_n272_), .C2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI22_X1  g079(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n268_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n264_), .A2(new_n282_), .A3(new_n276_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n266_), .B1(new_n283_), .B2(new_n267_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n265_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n232_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT34), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT35), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(KEYINPUT35), .ZN(new_n290_));
  AND4_X1   g089(.A1(new_n256_), .A2(new_n253_), .A3(new_n261_), .A4(new_n264_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n267_), .B1(new_n272_), .B2(new_n278_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT8), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n293_), .B2(new_n279_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n228_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .A4(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT35), .B(new_n288_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G218gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G134gat), .B(G162gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT73), .B(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT36), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n299_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(new_n299_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(KEYINPUT36), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n314_), .A2(KEYINPUT75), .A3(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n307_), .B(new_n313_), .C1(new_n316_), .C2(new_n312_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G64gat), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n320_));
  XOR2_X1   g119(.A(G71gat), .B(G78gat), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n222_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G231gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G183gat), .B(G211gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(KEYINPUT17), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(KEYINPUT17), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n327_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n333_), .B2(new_n327_), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT78), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n311_), .A2(new_n307_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n315_), .B1(new_n338_), .B2(KEYINPUT75), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n317_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT79), .Z(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  OAI22_X1  g141(.A1(new_n294_), .A2(new_n324_), .B1(KEYINPUT67), .B2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(KEYINPUT67), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n294_), .B2(new_n324_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n324_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n342_), .A2(KEYINPUT67), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n285_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT66), .B1(new_n285_), .B2(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n285_), .A2(new_n346_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  OAI21_X1  g152(.A(new_n350_), .B1(new_n353_), .B2(new_n349_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G176gat), .B(G204gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G120gat), .B(G148gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n354_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT13), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n341_), .A2(KEYINPUT80), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT90), .B(G197gat), .ZN(new_n366_));
  INV_X1    g165(.A(G204gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(G197gat), .B2(new_n367_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(KEYINPUT92), .B2(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(KEYINPUT21), .B(new_n375_), .C1(new_n366_), .C2(G204gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT91), .Z(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n372_), .A2(new_n373_), .A3(new_n378_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT85), .B1(new_n382_), .B2(KEYINPUT23), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(KEYINPUT23), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(KEYINPUT85), .ZN(new_n385_));
  NOR3_X1   g184(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G169gat), .B(G176gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G190gat), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n388_), .A2(KEYINPUT24), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT84), .B(G176gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n393_), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n384_), .B1(G183gat), .B2(G190gat), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n387_), .A2(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n381_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n386_), .B1(new_n391_), .B2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n384_), .C1(new_n399_), .C2(new_n391_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n385_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n381_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n397_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n381_), .A2(new_n396_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n379_), .A2(new_n380_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n404_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n412_), .A4(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT18), .B(G64gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  AND3_X1   g218(.A1(new_n410_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n365_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT102), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT102), .B(new_n365_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n419_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT101), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n411_), .A2(new_n414_), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n430_));
  OAI21_X1  g229(.A(new_n409_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n397_), .A2(new_n406_), .A3(KEYINPUT101), .A4(new_n412_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n420_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n424_), .A2(new_n425_), .B1(KEYINPUT27), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G127gat), .B(G134gat), .ZN(new_n436_));
  INV_X1    g235(.A(G113gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G120gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G155gat), .B(G162gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(KEYINPUT88), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(KEYINPUT88), .ZN(new_n442_));
  OR3_X1    g241(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444_));
  INV_X1    g243(.A(G141gat), .ZN(new_n445_));
  INV_X1    g244(.A(G148gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n442_), .A3(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n452_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n453_));
  OAI221_X1 g252(.A(new_n453_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n439_), .B2(new_n455_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n457_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n456_), .A2(KEYINPUT4), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT96), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT96), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n460_), .B2(KEYINPUT4), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n466_), .B2(new_n463_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n462_), .B1(new_n467_), .B2(new_n461_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G1gat), .B(G29gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G85gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n462_), .B(new_n475_), .C1(new_n467_), .C2(new_n461_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G228gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT89), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n455_), .A2(KEYINPUT29), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n413_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G78gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(new_n455_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n413_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  OAI21_X1  g290(.A(G78gat), .B1(new_n491_), .B2(new_n484_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(G106gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(G106gat), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n479_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n493_), .A3(KEYINPUT94), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n455_), .A2(KEYINPUT29), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(new_n227_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT28), .B(G22gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n404_), .B(new_n251_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT30), .Z(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G71gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n507_), .B(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n504_), .A2(new_n510_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n439_), .B(KEYINPUT31), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n513_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n502_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n479_), .B(new_n520_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n503_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n503_), .B2(new_n521_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n435_), .B(new_n478_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n503_), .A2(new_n521_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n433_), .A2(KEYINPUT32), .A3(new_n419_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT98), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n410_), .A2(new_n415_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n477_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n461_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n460_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n473_), .B(new_n534_), .C1(new_n467_), .C2(new_n533_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n410_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n410_), .A2(new_n415_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n426_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n476_), .A2(KEYINPUT33), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n476_), .A2(KEYINPUT33), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n519_), .B(new_n525_), .C1(new_n532_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n524_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n341_), .A2(new_n363_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AND4_X1   g346(.A1(new_n247_), .A2(new_n364_), .A3(new_n544_), .A4(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n211_), .A3(new_n477_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n363_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(new_n246_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n337_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n338_), .B(KEYINPUT103), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n544_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G1gat), .B1(new_n558_), .B2(new_n478_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n549_), .A2(new_n550_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n559_), .A3(new_n560_), .ZN(G1324gat));
  INV_X1    g360(.A(new_n435_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n548_), .A2(new_n212_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n564_));
  OAI211_X1 g363(.A(G8gat), .B(new_n564_), .C1(new_n558_), .C2(new_n435_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(G1325gat));
  INV_X1    g370(.A(G15gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n519_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n548_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n557_), .B2(new_n573_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT41), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(G1326gat));
  INV_X1    g376(.A(G22gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n525_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n557_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT42), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n548_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(G1327gat));
  AOI21_X1  g382(.A(new_n338_), .B1(new_n524_), .B2(new_n543_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n552_), .A2(new_n246_), .A3(new_n337_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(G29gat), .B1(new_n586_), .B2(new_n477_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT43), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n317_), .A2(new_n339_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT105), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n544_), .B2(new_n589_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n589_), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n594_), .B(new_n591_), .C1(new_n524_), .C2(new_n543_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(KEYINPUT44), .A3(new_n585_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n597_), .A2(new_n477_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n585_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT44), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(G29gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n587_), .B1(new_n598_), .B2(new_n602_), .ZN(G1328gat));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n562_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G36gat), .ZN(new_n605_));
  INV_X1    g404(.A(G36gat), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n562_), .A2(KEYINPUT106), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n562_), .A2(KEYINPUT106), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n586_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT45), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n605_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n605_), .B(new_n612_), .C1(KEYINPUT107), .C2(KEYINPUT46), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1329gat));
  NAND2_X1  g416(.A1(new_n597_), .A2(new_n573_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n601_), .A2(G43gat), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n586_), .A2(new_n573_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n618_), .A2(new_n619_), .B1(G43gat), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g421(.A(G50gat), .B1(new_n586_), .B2(new_n579_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n597_), .A2(new_n579_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n227_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n624_), .B2(new_n625_), .ZN(G1331gat));
  NOR2_X1   g425(.A1(new_n363_), .A2(new_n247_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n544_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n341_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G57gat), .B1(new_n630_), .B2(new_n477_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT108), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n632_), .A3(new_n556_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n544_), .A2(new_n556_), .A3(new_n627_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT108), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n478_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n631_), .B1(new_n637_), .B2(G57gat), .ZN(G1332gat));
  OR3_X1    g437(.A1(new_n629_), .A2(G64gat), .A3(new_n609_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G64gat), .B1(new_n636_), .B2(new_n609_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT48), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(KEYINPUT48), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(G1333gat));
  NOR2_X1   g442(.A1(new_n519_), .A2(G71gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT109), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n630_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n573_), .A3(new_n635_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT49), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G71gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G71gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT110), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1334gat));
  NAND3_X1  g452(.A1(new_n630_), .A2(new_n486_), .A3(new_n579_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT50), .ZN(new_n655_));
  INV_X1    g454(.A(new_n636_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n579_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n657_), .B2(G78gat), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT50), .B(new_n486_), .C1(new_n656_), .C2(new_n579_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(G1335gat));
  NOR3_X1   g459(.A1(new_n363_), .A2(new_n247_), .A3(new_n337_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n584_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n257_), .B1(new_n662_), .B2(new_n478_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT111), .Z(new_n664_));
  AND2_X1   g463(.A1(new_n596_), .A2(new_n661_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n478_), .A2(new_n257_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(G1336gat));
  NAND3_X1  g466(.A1(new_n665_), .A2(G92gat), .A3(new_n610_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n258_), .B1(new_n662_), .B2(new_n435_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT112), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1337gat));
  NAND2_X1  g471(.A1(new_n596_), .A2(new_n661_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G99gat), .B1(new_n673_), .B2(new_n519_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n573_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n662_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g476(.A(new_n579_), .B(new_n661_), .C1(new_n593_), .C2(new_n595_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G106gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT113), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT113), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n681_), .A3(G106gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n680_), .A2(KEYINPUT52), .A3(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n584_), .A2(new_n248_), .A3(new_n579_), .A4(new_n661_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT52), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(KEYINPUT113), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT53), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT53), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n683_), .A2(new_n689_), .A3(new_n684_), .A4(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1339gat));
  INV_X1    g490(.A(KEYINPUT114), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n350_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT55), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n343_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n349_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT115), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT55), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n350_), .A2(new_n692_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT115), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n701_), .A3(new_n696_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n694_), .A2(new_n698_), .A3(new_n700_), .A4(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n361_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT56), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n703_), .A2(KEYINPUT56), .A3(new_n361_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(KEYINPUT116), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT116), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n703_), .A2(new_n709_), .A3(KEYINPUT56), .A4(new_n361_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n354_), .A2(new_n361_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n712_), .A3(new_n247_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT117), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n234_), .A2(new_n235_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n225_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n206_), .B(new_n717_), .C1(new_n241_), .C2(new_n225_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n242_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n362_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n708_), .A2(new_n712_), .A3(new_n247_), .A4(KEYINPUT117), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n715_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n338_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT57), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(KEYINPUT57), .A3(new_n338_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n706_), .A2(new_n707_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n711_), .A3(new_n719_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT58), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n589_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n726_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n554_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n340_), .A2(new_n733_), .A3(new_n246_), .A4(new_n363_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n317_), .A2(new_n246_), .A3(new_n337_), .A4(new_n339_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT54), .B1(new_n735_), .B2(new_n552_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n435_), .A2(new_n525_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n478_), .A2(new_n519_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT59), .B1(new_n742_), .B2(KEYINPUT118), .ZN(new_n743_));
  OR2_X1    g542(.A1(KEYINPUT119), .A2(G113gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(G113gat), .B1(new_n246_), .B2(KEYINPUT119), .ZN(new_n745_));
  NOR2_X1   g544(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n738_), .A2(new_n740_), .A3(new_n741_), .A4(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n437_), .B1(new_n742_), .B2(new_n246_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1340gat));
  NAND3_X1  g549(.A1(new_n743_), .A2(new_n552_), .A3(new_n747_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT120), .B(G120gat), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT60), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n742_), .B1(new_n754_), .B2(new_n752_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n363_), .A2(KEYINPUT60), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n752_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(G1341gat));
  NAND4_X1  g557(.A1(new_n743_), .A2(G127gat), .A3(new_n337_), .A4(new_n747_), .ZN(new_n759_));
  INV_X1    g558(.A(G127gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n742_), .B2(new_n554_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1342gat));
  INV_X1    g561(.A(KEYINPUT121), .ZN(new_n763_));
  INV_X1    g562(.A(new_n737_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n731_), .B2(new_n554_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n741_), .ZN(new_n766_));
  NOR4_X1   g565(.A1(new_n765_), .A2(KEYINPUT118), .A3(new_n739_), .A4(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT59), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n589_), .B(new_n747_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G134gat), .ZN(new_n770_));
  INV_X1    g569(.A(G134gat), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n738_), .A2(new_n771_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n555_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n763_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT121), .B(new_n774_), .C1(new_n769_), .C2(G134gat), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1343gat));
  INV_X1    g577(.A(new_n522_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n765_), .A2(new_n478_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n609_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n247_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT122), .B(G141gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(G1344gat));
  NOR2_X1   g584(.A1(new_n781_), .A2(new_n363_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(new_n446_), .ZN(G1345gat));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n337_), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT61), .B(G155gat), .Z(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT123), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n788_), .B(new_n790_), .ZN(G1346gat));
  AOI21_X1  g590(.A(G162gat), .B1(new_n782_), .B2(new_n555_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n781_), .A2(new_n594_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(G162gat), .B2(new_n793_), .ZN(G1347gat));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n765_), .A2(new_n519_), .A3(new_n579_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n609_), .A2(new_n477_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n246_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n799_), .B2(new_n203_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n393_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT62), .B(G169gat), .C1(new_n798_), .C2(new_n246_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(G1348gat));
  AND2_X1   g602(.A1(new_n796_), .A2(new_n797_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(G176gat), .A3(new_n552_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n392_), .B1(new_n798_), .B2(new_n363_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT124), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n805_), .ZN(G1349gat));
  NOR2_X1   g609(.A1(new_n798_), .A2(new_n554_), .ZN(new_n811_));
  MUX2_X1   g610(.A(G183gat), .B(new_n389_), .S(new_n811_), .Z(G1350gat));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n390_), .A3(new_n555_), .ZN(new_n813_));
  OAI21_X1  g612(.A(G190gat), .B1(new_n798_), .B2(new_n594_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1351gat));
  NOR2_X1   g614(.A1(new_n765_), .A2(new_n779_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n797_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT125), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n819_), .A3(new_n797_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n246_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT126), .A3(new_n205_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT126), .B(G197gat), .Z(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(new_n823_), .ZN(G1352gat));
  NAND2_X1  g623(.A1(new_n818_), .A2(new_n820_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n552_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT127), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n367_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n825_), .A2(new_n552_), .B1(new_n827_), .B2(new_n367_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1353gat));
  XNOR2_X1  g630(.A(KEYINPUT63), .B(G211gat), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n554_), .B(new_n832_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n337_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1354gat));
  AOI21_X1  g635(.A(G218gat), .B1(new_n825_), .B2(new_n555_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n594_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(G218gat), .B2(new_n838_), .ZN(G1355gat));
endmodule


