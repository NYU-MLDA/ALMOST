//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(G57gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G64gat), .ZN(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G57gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(G57gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(G64gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT64), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n202_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n202_), .A3(new_n211_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G71gat), .B(G78gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n215_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT64), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n209_), .B2(new_n210_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT65), .B1(new_n223_), .B2(new_n216_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n212_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G231gat), .A3(G233gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G231gat), .A2(G233gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G8gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT75), .ZN(new_n233_));
  INV_X1    g032(.A(G15gat), .ZN(new_n234_));
  INV_X1    g033(.A(G22gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G15gat), .A2(G22gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G1gat), .A2(G8gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n236_), .A2(new_n237_), .B1(KEYINPUT14), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n233_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n231_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n240_), .A3(new_n230_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G127gat), .B(G155gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(G183gat), .B(G211gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT77), .B1(new_n242_), .B2(new_n244_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n243_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G29gat), .B(G36gat), .Z(new_n261_));
  XOR2_X1   g060(.A(G43gat), .B(G50gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT79), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(new_n241_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G229gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n263_), .B(KEYINPUT15), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n240_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n264_), .B2(new_n241_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n265_), .A2(new_n267_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G113gat), .B(G141gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(G169gat), .B(G197gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n271_), .B(new_n274_), .Z(new_n275_));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT81), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT24), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n279_), .A2(KEYINPUT24), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT23), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  INV_X1    g086(.A(G190gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT80), .B1(new_n288_), .B2(KEYINPUT26), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n287_), .B(new_n289_), .C1(new_n290_), .C2(KEYINPUT80), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n281_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT22), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(KEYINPUT22), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n293_), .B(new_n296_), .C1(new_n297_), .C2(new_n294_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT83), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT84), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n285_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n283_), .A2(new_n285_), .A3(new_n300_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n279_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n292_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT30), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT85), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G71gat), .B(G99gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G43gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(new_n234_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n310_), .B(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n307_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n318_), .A2(KEYINPUT86), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(KEYINPUT86), .ZN(new_n320_));
  XOR2_X1   g119(.A(G113gat), .B(G120gat), .Z(new_n321_));
  OR3_X1    g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n314_), .A2(new_n317_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G141gat), .ZN(new_n334_));
  INV_X1    g133(.A(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n333_), .A2(KEYINPUT2), .B1(new_n336_), .B2(KEYINPUT3), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(KEYINPUT88), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OAI221_X1 g140(.A(new_n337_), .B1(KEYINPUT3), .B2(new_n336_), .C1(KEYINPUT2), .C2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G155gat), .B(G162gat), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n336_), .B(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n341_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT29), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT28), .Z(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  XOR2_X1   g154(.A(G197gat), .B(G204gat), .Z(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT21), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(KEYINPUT21), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n358_), .A2(new_n359_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n351_), .A2(KEYINPUT29), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n366_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n355_), .A2(KEYINPUT90), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(KEYINPUT90), .B2(new_n355_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n355_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n367_), .A2(KEYINPUT91), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(KEYINPUT91), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .A4(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n351_), .B(new_n324_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT4), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT99), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n351_), .A2(new_n324_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT4), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n377_), .B(new_n379_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n378_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n385_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n360_), .A2(new_n361_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n306_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n290_), .A2(new_n287_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n281_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n304_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT93), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT22), .B(G169gat), .Z(new_n406_));
  OAI21_X1  g205(.A(new_n279_), .B1(new_n406_), .B2(G176gat), .ZN(new_n407_));
  OAI22_X1  g206(.A1(new_n403_), .A2(new_n303_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n408_), .B2(new_n399_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n401_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n408_), .B2(new_n399_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n399_), .B2(new_n306_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n398_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT96), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(KEYINPUT32), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n413_), .A2(new_n398_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT94), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n408_), .A2(new_n423_), .A3(new_n399_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n408_), .B2(new_n399_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n398_), .A2(new_n411_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .A4(new_n400_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n395_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n377_), .B(new_n378_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n376_), .A2(new_n379_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n393_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n391_), .A2(KEYINPUT33), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n386_), .A2(new_n437_), .A3(new_n390_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n422_), .A2(new_n427_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n420_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n422_), .A2(new_n427_), .A3(new_n420_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT97), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n445_), .A3(new_n441_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(KEYINPUT98), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT98), .B1(new_n444_), .B2(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n439_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n431_), .B1(new_n450_), .B2(KEYINPUT101), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n437_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n392_), .A2(KEYINPUT33), .A3(new_n393_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n434_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n444_), .A2(new_n446_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT98), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n447_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT101), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n375_), .B1(new_n451_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n395_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n375_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n444_), .A2(new_n464_), .A3(new_n446_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n414_), .A2(new_n441_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT27), .A3(new_n443_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n331_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n395_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n370_), .A2(new_n374_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT102), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT102), .B1(new_n465_), .B2(new_n467_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n471_), .B(new_n472_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT103), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n275_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G230gat), .A2(G233gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n482_), .A2(KEYINPUT9), .ZN(new_n483_));
  OR2_X1    g282(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(KEYINPUT9), .A3(new_n482_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n481_), .A2(new_n483_), .A3(new_n487_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n490_), .A2(new_n482_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n480_), .B(new_n495_), .ZN(new_n496_));
  OR3_X1    g295(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n494_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n493_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n220_), .A2(new_n226_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n504_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n218_), .A2(new_n219_), .A3(new_n213_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n212_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n479_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n504_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT68), .B1(new_n513_), .B2(KEYINPUT12), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT12), .B(new_n508_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(KEYINPUT67), .A3(KEYINPUT12), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n514_), .A2(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n505_), .A2(new_n479_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n512_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G120gat), .B(G148gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n524_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n268_), .A2(new_n508_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n504_), .A2(new_n263_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n540_), .B1(KEYINPUT35), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n537_), .B2(KEYINPUT71), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT72), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT73), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n554_), .B(new_n555_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT74), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n550_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n548_), .A2(KEYINPUT74), .A3(new_n549_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n550_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(KEYINPUT37), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n564_), .A2(KEYINPUT37), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND4_X1   g367(.A1(new_n260_), .A2(new_n478_), .A3(new_n536_), .A4(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G1gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n395_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT38), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n564_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n535_), .A2(new_n259_), .A3(new_n275_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT104), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT104), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n577_), .A3(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n462_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n572_), .A2(new_n581_), .ZN(G1324gat));
  INV_X1    g381(.A(G8gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n473_), .A2(new_n474_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n569_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G8gat), .B1(new_n575_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g390(.A(new_n234_), .B1(new_n579_), .B2(new_n330_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n569_), .A2(new_n234_), .A3(new_n330_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(G1326gat));
  NAND3_X1  g396(.A1(new_n569_), .A2(new_n235_), .A3(new_n375_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G22gat), .B1(new_n580_), .B2(new_n472_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT42), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(KEYINPUT42), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(G1327gat));
  AOI21_X1  g401(.A(new_n568_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT43), .B1(new_n603_), .B2(KEYINPUT106), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n430_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n450_), .A2(KEYINPUT101), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n472_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n469_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n330_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n475_), .B(KEYINPUT103), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n567_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n535_), .A2(new_n275_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n604_), .A2(new_n614_), .A3(new_n259_), .A4(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n611_), .A2(new_n612_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n260_), .B1(new_n619_), .B2(KEYINPUT43), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(KEYINPUT44), .A3(new_n615_), .A4(new_n614_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n618_), .A2(new_n621_), .A3(G29gat), .A4(new_n395_), .ZN(new_n622_));
  INV_X1    g421(.A(G29gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n564_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n260_), .A2(new_n535_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n478_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT108), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n478_), .A2(KEYINPUT108), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n623_), .B1(new_n630_), .B2(new_n462_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n622_), .A2(new_n631_), .ZN(G1328gat));
  NAND3_X1  g431(.A1(new_n618_), .A2(new_n621_), .A3(new_n584_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n586_), .A2(G36gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT45), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT46), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(KEYINPUT46), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n618_), .A2(new_n621_), .A3(G43gat), .A4(new_n330_), .ZN(new_n643_));
  INV_X1    g442(.A(G43gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n630_), .B2(new_n331_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g446(.A1(new_n618_), .A2(new_n621_), .A3(G50gat), .A4(new_n375_), .ZN(new_n648_));
  INV_X1    g447(.A(G50gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n630_), .B2(new_n472_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1331gat));
  INV_X1    g450(.A(new_n275_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n260_), .A2(new_n653_), .A3(new_n535_), .A4(new_n568_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n204_), .A3(new_n395_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n260_), .A2(new_n275_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n536_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n573_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n573_), .A2(KEYINPUT109), .A3(new_n657_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n395_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n662_), .B2(new_n204_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT110), .Z(G1332gat));
  NAND3_X1  g463(.A1(new_n654_), .A2(new_n206_), .A3(new_n584_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n584_), .A3(new_n661_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT48), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G64gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G64gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1333gat));
  INV_X1    g469(.A(G71gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n654_), .A2(new_n671_), .A3(new_n330_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n660_), .A2(new_n330_), .A3(new_n661_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT49), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(G71gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n673_), .B2(G71gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT111), .ZN(G1334gat));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n654_), .A2(new_n679_), .A3(new_n375_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n660_), .A2(new_n375_), .A3(new_n661_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT50), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G78gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G78gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1335gat));
  NOR2_X1   g484(.A1(new_n536_), .A2(new_n652_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n604_), .A2(new_n614_), .A3(new_n259_), .A4(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G85gat), .B1(new_n687_), .B2(new_n462_), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n564_), .A2(new_n653_), .A3(new_n259_), .A4(new_n535_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n488_), .A3(new_n395_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1336gat));
  OAI21_X1  g490(.A(G92gat), .B1(new_n687_), .B2(new_n586_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n489_), .A3(new_n584_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1337gat));
  NAND4_X1  g493(.A1(new_n689_), .A2(new_n330_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT112), .B(G99gat), .C1(new_n687_), .C2(new_n331_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n620_), .A2(new_n330_), .A3(new_n614_), .A4(new_n686_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT112), .B1(new_n698_), .B2(G99gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT51), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n695_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n689_), .A2(new_n485_), .A3(new_n375_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n485_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n706_), .B(new_n707_), .C1(new_n687_), .C2(new_n472_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n620_), .A2(new_n375_), .A3(new_n614_), .A4(new_n686_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n705_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT53), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n705_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1339gat));
  NOR2_X1   g515(.A1(new_n567_), .A2(new_n535_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n656_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n260_), .A2(KEYINPUT114), .A3(new_n275_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .A4(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n524_), .A2(new_n530_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n275_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n517_), .A2(new_n514_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n520_), .A2(new_n521_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n523_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n737_));
  NAND2_X1  g536(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n479_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n522_), .B2(new_n507_), .ZN(new_n743_));
  AND4_X1   g542(.A1(new_n742_), .A2(new_n730_), .A3(new_n731_), .A4(new_n507_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n729_), .B(new_n530_), .C1(new_n740_), .C2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n732_), .A2(new_n738_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n737_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n749_), .A3(new_n735_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n529_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n728_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n271_), .A2(new_n274_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n274_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n264_), .A2(new_n241_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n269_), .A3(new_n267_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n531_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n564_), .B1(new_n752_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT57), .B1(new_n761_), .B2(KEYINPUT118), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n749_), .A2(new_n735_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n730_), .A2(new_n731_), .A3(new_n507_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT117), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n522_), .A2(new_n742_), .A3(new_n507_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n479_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n529_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n729_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n529_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n773_), .A2(new_n728_), .B1(new_n531_), .B2(new_n759_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n763_), .B(new_n764_), .C1(new_n774_), .C2(new_n564_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n727_), .A2(new_n758_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(KEYINPUT58), .A3(new_n776_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n567_), .A3(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n762_), .A2(new_n775_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n260_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n762_), .A2(new_n775_), .A3(KEYINPUT119), .A4(new_n781_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n726_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n584_), .A2(new_n375_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n395_), .A3(new_n330_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT59), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n782_), .A2(new_n259_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n726_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n782_), .A2(new_n783_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n259_), .A3(new_n785_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n726_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n788_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT59), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT121), .B(new_n792_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n795_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(G113gat), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n275_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G113gat), .B1(new_n799_), .B2(new_n652_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT120), .Z(new_n806_));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1340gat));
  INV_X1    g606(.A(G120gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n536_), .B2(KEYINPUT60), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n799_), .B(new_n809_), .C1(KEYINPUT60), .C2(new_n808_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n789_), .A2(new_n535_), .A3(new_n792_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(new_n808_), .ZN(G1341gat));
  OAI21_X1  g612(.A(G127gat), .B1(new_n802_), .B2(new_n259_), .ZN(new_n814_));
  INV_X1    g613(.A(G127gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n799_), .A2(new_n815_), .A3(new_n260_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1342gat));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n818_));
  INV_X1    g617(.A(new_n801_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n789_), .B2(new_n792_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n567_), .A2(G134gat), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G134gat), .B1(new_n799_), .B2(new_n564_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT122), .B(new_n825_), .C1(new_n802_), .C2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1343gat));
  NOR2_X1   g626(.A1(new_n786_), .A2(new_n330_), .ZN(new_n828_));
  AND4_X1   g627(.A1(new_n395_), .A2(new_n828_), .A3(new_n375_), .A4(new_n586_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n652_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n535_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n260_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT61), .B(G155gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1346gat));
  AOI21_X1  g635(.A(G162gat), .B1(new_n829_), .B2(new_n564_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n567_), .A2(G162gat), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT123), .Z(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n829_), .B2(new_n839_), .ZN(G1347gat));
  NOR2_X1   g639(.A1(new_n791_), .A2(new_n726_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n584_), .A2(new_n471_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n472_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n846_), .A2(new_n406_), .A3(new_n275_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n295_), .B1(new_n845_), .B2(new_n652_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(KEYINPUT62), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(KEYINPUT62), .B2(new_n848_), .ZN(G1348gat));
  AOI21_X1  g649(.A(G176gat), .B1(new_n845_), .B2(new_n535_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n786_), .A2(new_n375_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n843_), .A2(G176gat), .A3(new_n535_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  NOR3_X1   g653(.A1(new_n846_), .A2(new_n287_), .A3(new_n259_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n852_), .A2(new_n260_), .A3(new_n843_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT125), .ZN(new_n857_));
  AOI21_X1  g656(.A(G183gat), .B1(new_n856_), .B2(KEYINPUT125), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n846_), .B2(new_n568_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n845_), .A2(new_n290_), .A3(new_n564_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1351gat));
  NOR2_X1   g661(.A1(new_n586_), .A2(new_n463_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n828_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n652_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n535_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g668(.A1(new_n864_), .A2(new_n259_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n870_), .A2(KEYINPUT126), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT126), .B1(new_n870_), .B2(new_n872_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT63), .B(G211gat), .Z(new_n875_));
  AOI22_X1  g674(.A1(new_n873_), .A2(new_n874_), .B1(new_n870_), .B2(new_n875_), .ZN(G1354gat));
  OR3_X1    g675(.A1(new_n864_), .A2(G218gat), .A3(new_n624_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G218gat), .B1(new_n864_), .B2(new_n568_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1355gat));
endmodule


