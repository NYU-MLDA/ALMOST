//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT85), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n202_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT84), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n206_), .A2(new_n207_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT86), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n207_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(G169gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G183gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n203_), .A2(new_n205_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n230_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT24), .A3(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n220_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(KEYINPUT88), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G15gat), .B(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT87), .ZN(new_n241_));
  INV_X1    g040(.A(G99gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G71gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n238_), .B2(KEYINPUT88), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n239_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250_));
  INV_X1    g049(.A(G120gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G113gat), .ZN(new_n252_));
  INV_X1    g051(.A(G113gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G120gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G134gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G127gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G134gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT90), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT90), .B1(new_n257_), .B2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n255_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n258_), .A2(G134gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n256_), .A2(G127gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT90), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n252_), .A2(new_n254_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n250_), .B1(new_n271_), .B2(KEYINPUT89), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n250_), .B2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n249_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n239_), .A2(new_n248_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n239_), .A2(new_n248_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G197gat), .A2(G204gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(KEYINPUT21), .A3(new_n280_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT93), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n293_), .A2(new_n294_), .B1(new_n289_), .B2(KEYINPUT1), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT93), .A3(G155gat), .A4(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(KEYINPUT92), .A3(KEYINPUT1), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n292_), .A2(new_n295_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300_));
  OR3_X1    g099(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  INV_X1    g101(.A(G141gat), .ZN(new_n303_));
  INV_X1    g102(.A(G148gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n301_), .A2(new_n305_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n293_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(new_n289_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n299_), .A2(new_n300_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n288_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G228gat), .ZN(new_n314_));
  INV_X1    g113(.A(G233gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  OAI221_X1 g116(.A(new_n288_), .B1(new_n314_), .B2(new_n315_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G78gat), .B(G106gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT95), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n311_), .A2(new_n312_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G22gat), .B(G50gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n323_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n320_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n317_), .A2(new_n318_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n322_), .A2(new_n321_), .A3(new_n330_), .A4(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT99), .B1(new_n311_), .B2(new_n270_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n299_), .A2(new_n300_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n308_), .A2(new_n310_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n260_), .A2(new_n261_), .A3(new_n255_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n268_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n342_), .A3(KEYINPUT99), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G85gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT0), .B(G57gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  INV_X1    g151(.A(new_n347_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n311_), .A2(new_n270_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT100), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT100), .ZN(new_n357_));
  NOR4_X1   g156(.A1(new_n311_), .A2(new_n270_), .A3(new_n357_), .A4(KEYINPUT4), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n355_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n348_), .B(new_n352_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT33), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n346_), .A2(KEYINPUT4), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n357_), .B1(new_n343_), .B2(KEYINPUT4), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n354_), .A2(KEYINPUT100), .A3(new_n355_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n347_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n348_), .A4(new_n352_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G8gat), .B(G36gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT18), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n286_), .A2(new_n287_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n220_), .B2(new_n236_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT19), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n212_), .A2(new_n208_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n229_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n219_), .ZN(new_n381_));
  AND2_X1   g180(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n221_), .B(new_n223_), .C1(new_n382_), .C2(new_n227_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n231_), .A2(KEYINPUT96), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT24), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n386_), .A3(new_n230_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n233_), .A2(new_n234_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n383_), .B(new_n387_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n206_), .A2(new_n207_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n381_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT20), .B(new_n378_), .C1(new_n392_), .C2(new_n288_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n220_), .A2(new_n236_), .A3(new_n375_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n392_), .B2(new_n288_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n378_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n394_), .A2(new_n395_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT97), .B1(new_n376_), .B2(new_n393_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n374_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n393_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n237_), .A2(new_n288_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n400_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n374_), .A2(new_n406_), .A3(new_n402_), .A4(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT98), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(new_n374_), .A3(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n374_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n352_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n347_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n360_), .B2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n370_), .A2(new_n409_), .A3(new_n415_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n367_), .A2(new_n348_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n352_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n361_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n288_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n400_), .B1(new_n376_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n396_), .A2(new_n398_), .A3(new_n378_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n374_), .A2(KEYINPUT32), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n411_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n411_), .B2(KEYINPUT101), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n335_), .B1(new_n419_), .B2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n422_), .A2(new_n332_), .A3(new_n333_), .A4(new_n361_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n374_), .B(KEYINPUT102), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n410_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n278_), .B1(new_n435_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT103), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n278_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n423_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n335_), .A2(new_n442_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT103), .B(new_n278_), .C1(new_n435_), .C2(new_n443_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G229gat), .A2(G233gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT71), .B(G1gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(G8gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(G15gat), .B(G22gat), .Z(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT72), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(G8gat), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT14), .ZN(new_n464_));
  INV_X1    g263(.A(new_n459_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n460_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G36gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G29gat), .ZN(new_n474_));
  INV_X1    g273(.A(G29gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(G36gat), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n474_), .A2(new_n476_), .A3(KEYINPUT69), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT69), .B1(new_n474_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n472_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n476_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n474_), .A2(new_n476_), .A3(KEYINPUT69), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n471_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n469_), .A2(new_n470_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n468_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n458_), .A2(KEYINPUT72), .A3(new_n459_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n466_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n460_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n455_), .B1(new_n486_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n485_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT77), .A3(new_n455_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n479_), .A2(new_n484_), .A3(KEYINPUT15), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT15), .B1(new_n479_), .B2(new_n484_), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n469_), .A2(new_n470_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n499_), .A3(new_n454_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n504_), .A2(KEYINPUT78), .A3(new_n499_), .A4(new_n454_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n496_), .A2(new_n501_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT79), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G113gat), .B(G141gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT80), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT81), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n453_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n509_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n496_), .A2(new_n501_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n507_), .A2(new_n508_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT79), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n526_), .A2(new_n511_), .A3(KEYINPUT82), .A4(new_n518_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT83), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n520_), .A2(new_n530_), .A3(new_n522_), .A4(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n452_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(G183gat), .B(G211gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT17), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n497_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n497_), .A2(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT73), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n539_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(KEYINPUT74), .A3(new_n556_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT74), .ZN(new_n559_));
  INV_X1    g358(.A(new_n550_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n552_), .B1(new_n560_), .B2(new_n548_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT76), .Z(new_n565_));
  AOI21_X1  g364(.A(new_n557_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT10), .B(G99gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G106gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(KEYINPUT65), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n571_));
  INV_X1    g370(.A(G85gat), .ZN(new_n572_));
  INV_X1    g371(.A(G92gat), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(G85gat), .B(G92gat), .C1(KEYINPUT66), .C2(KEYINPUT9), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT6), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(G99gat), .A3(G106gat), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n574_), .A2(new_n575_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT65), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n567_), .B2(G106gat), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n570_), .A2(new_n576_), .A3(new_n581_), .A4(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n580_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(new_n242_), .A3(new_n569_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT8), .ZN(new_n590_));
  XOR2_X1   g389(.A(G85gat), .B(G92gat), .Z(new_n591_));
  AND3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n584_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n547_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n546_), .B(new_n584_), .C1(new_n593_), .C2(new_n592_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT12), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n547_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT64), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G176gat), .B(G204gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT68), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n604_), .A2(new_n606_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT13), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n566_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n622_));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n594_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT34), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n487_), .B(new_n584_), .C1(new_n593_), .C2(new_n592_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n629_), .A2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n626_), .A2(new_n636_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n622_), .B(new_n625_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT70), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n625_), .A2(new_n622_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n638_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n644_), .A2(new_n645_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n621_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n533_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(new_n448_), .A3(new_n457_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT38), .Z(new_n651_));
  AND2_X1   g450(.A1(new_n452_), .A2(new_n644_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n528_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n618_), .A2(new_n620_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n657_), .B2(new_n528_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n566_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n652_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n423_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G1gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n651_), .A2(new_n666_), .ZN(G1324gat));
  NAND3_X1  g466(.A1(new_n652_), .A2(new_n660_), .A3(new_n442_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n671_), .A3(G8gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n672_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n442_), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n649_), .A2(G8gat), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n675_), .A2(new_n677_), .A3(new_n679_), .A4(new_n681_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  OR3_X1    g484(.A1(new_n649_), .A2(G15gat), .A3(new_n278_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n663_), .A2(new_n447_), .A3(new_n664_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n687_), .B2(G15gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1326gat));
  OR3_X1    g489(.A1(new_n649_), .A2(G22gat), .A3(new_n334_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n663_), .A2(new_n335_), .A3(new_n664_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G22gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G22gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n644_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n657_), .A2(new_n697_), .A3(new_n659_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n533_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n423_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n646_), .A2(new_n647_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n419_), .A2(new_n434_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n334_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n443_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT103), .B1(new_n708_), .B2(new_n278_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n451_), .A2(new_n450_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n703_), .B(new_n704_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n452_), .A2(KEYINPUT109), .A3(new_n703_), .A4(new_n704_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n704_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT43), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n656_), .A2(new_n658_), .A3(new_n566_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n448_), .A2(new_n475_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n702_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n721_), .A2(new_n442_), .A3(new_n722_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n473_), .A2(KEYINPUT110), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n678_), .A2(G36gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n533_), .A2(new_n699_), .A3(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT45), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n731_), .B2(KEYINPUT45), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n726_), .B1(new_n729_), .B2(new_n736_), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT46), .B(new_n735_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  NAND4_X1  g538(.A1(new_n721_), .A2(G43gat), .A3(new_n447_), .A4(new_n722_), .ZN(new_n740_));
  INV_X1    g539(.A(G43gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n700_), .B2(new_n278_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT47), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n745_), .A3(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n701_), .B2(new_n335_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n335_), .A2(G50gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n723_), .B2(new_n749_), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n532_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n652_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n448_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n452_), .A2(new_n653_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n704_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n655_), .A3(new_n566_), .A4(new_n755_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n448_), .A2(G57gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1332gat));
  OAI21_X1  g557(.A(G64gat), .B1(new_n752_), .B2(new_n678_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n678_), .A2(G64gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n756_), .B2(new_n762_), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n752_), .B2(new_n278_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT49), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n447_), .A2(new_n245_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n756_), .B2(new_n766_), .ZN(G1334gat));
  OAI21_X1  g566(.A(G78gat), .B1(new_n752_), .B2(new_n334_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT50), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n334_), .A2(G78gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n756_), .B2(new_n770_), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n657_), .A2(new_n566_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n754_), .A2(new_n697_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n572_), .A3(new_n423_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n653_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT112), .Z(new_n777_));
  NAND2_X1  g576(.A1(new_n717_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n717_), .A2(KEYINPUT113), .A3(new_n777_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n448_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n775_), .B1(new_n782_), .B2(new_n572_), .ZN(G1336gat));
  OAI21_X1  g582(.A(new_n573_), .B1(new_n773_), .B2(new_n678_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT114), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n442_), .A2(G92gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT115), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n785_), .B1(new_n786_), .B2(new_n788_), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n774_), .A2(new_n447_), .A3(new_n568_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n278_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n242_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n790_), .C1(new_n791_), .C2(new_n242_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1338gat));
  OAI21_X1  g595(.A(G106gat), .B1(new_n778_), .B2(new_n334_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(G106gat), .B(new_n802_), .C1(new_n778_), .C2(new_n334_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n774_), .A2(new_n569_), .A3(new_n335_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n800_), .A2(new_n807_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n648_), .A2(new_n531_), .A3(new_n529_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n500_), .A2(new_n454_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n504_), .A2(new_n499_), .A3(new_n455_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n516_), .A3(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n522_), .A2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n818_), .A2(new_n617_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n597_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n602_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n600_), .A2(new_n823_), .A3(new_n603_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n614_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n820_), .B(KEYINPUT56), .C1(new_n824_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n616_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n597_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n604_), .A2(KEYINPUT55), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n613_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n820_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n828_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n819_), .B1(new_n528_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n814_), .B1(new_n835_), .B2(new_n697_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n522_), .A2(new_n616_), .A3(new_n817_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n522_), .A2(KEYINPUT119), .A3(new_n616_), .A4(new_n817_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n831_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n839_), .A2(new_n840_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT120), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(KEYINPUT120), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n839_), .A2(new_n848_), .A3(new_n840_), .A4(new_n844_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n704_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n527_), .A2(new_n522_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n517_), .B1(new_n525_), .B2(KEYINPUT79), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT82), .B1(new_n853_), .B2(new_n511_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n834_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n819_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n697_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n851_), .B1(new_n857_), .B2(KEYINPUT57), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n835_), .A2(KEYINPUT121), .A3(new_n814_), .A4(new_n697_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n836_), .B(new_n850_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n813_), .B1(new_n860_), .B2(new_n659_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n447_), .A2(new_n423_), .A3(new_n449_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n811_), .B(KEYINPUT54), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n850_), .B1(new_n857_), .B2(KEYINPUT57), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n855_), .A2(new_n856_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT121), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n857_), .A2(new_n851_), .A3(KEYINPUT57), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n865_), .B1(new_n871_), .B2(new_n566_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n863_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n810_), .B1(new_n864_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n862_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(KEYINPUT59), .A3(new_n873_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(KEYINPUT122), .A3(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n532_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G113gat), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n861_), .A2(new_n863_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n253_), .A3(new_n528_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1340gat));
  OAI21_X1  g682(.A(new_n251_), .B1(new_n657_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n881_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n251_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n657_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G120gat), .B1(new_n886_), .B2(new_n887_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1341gat));
  NAND3_X1  g689(.A1(new_n875_), .A2(new_n566_), .A3(new_n878_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G127gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n881_), .A2(new_n258_), .A3(new_n566_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1342gat));
  NAND3_X1  g693(.A1(new_n875_), .A2(new_n704_), .A3(new_n878_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G134gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n881_), .A2(new_n256_), .A3(new_n697_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1343gat));
  NOR3_X1   g697(.A1(new_n447_), .A2(new_n448_), .A3(new_n334_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n872_), .A2(new_n678_), .A3(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n653_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT124), .B(G141gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1344gat));
  NOR2_X1   g702(.A1(new_n900_), .A2(new_n657_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n304_), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n900_), .A2(new_n659_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT61), .B(G155gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n900_), .B2(new_n755_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n644_), .A2(G162gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n900_), .B2(new_n910_), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n861_), .A2(new_n678_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n278_), .A2(new_n423_), .A3(new_n335_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n528_), .A3(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n914_), .B2(KEYINPUT22), .ZN(new_n915_));
  OAI21_X1  g714(.A(G169gat), .B1(new_n914_), .B2(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(G169gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n915_), .ZN(G1348gat));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n913_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n657_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(G176gat), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(G176gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT125), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n921_), .B2(new_n925_), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n912_), .A2(new_n566_), .A3(new_n913_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n224_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n212_), .B2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n920_), .B2(new_n755_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n697_), .B1(new_n227_), .B2(new_n382_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n920_), .B2(new_n931_), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n447_), .A2(new_n436_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n912_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n528_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT126), .B(G197gat), .Z(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1352gat));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n655_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n912_), .A2(new_n566_), .A3(new_n933_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n940_), .B2(new_n941_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n934_), .B2(new_n697_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n704_), .A2(G218gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT127), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n934_), .B2(new_n947_), .ZN(G1355gat));
endmodule


