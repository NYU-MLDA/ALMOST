//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT25), .B(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT77), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT23), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n214_), .A2(new_n222_), .A3(KEYINPUT23), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n218_), .A2(new_n219_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n213_), .B1(new_n221_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n229_), .A3(new_n208_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(KEYINPUT79), .A3(new_n208_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n232_), .A2(new_n234_), .A3(new_n210_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n214_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n215_), .A2(new_n217_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n237_), .B(new_n239_), .C1(new_n241_), .C2(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT80), .ZN(new_n249_));
  XOR2_X1   g048(.A(G15gat), .B(G43gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(KEYINPUT81), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n246_), .A2(KEYINPUT82), .A3(new_n255_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT82), .B1(new_n246_), .B2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n262_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT31), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n257_), .A2(new_n260_), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n202_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n257_), .A2(new_n260_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n257_), .A2(new_n260_), .A3(new_n268_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT84), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G228gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G78gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G106gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G22gat), .B(G50gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT3), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT2), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n290_), .B2(KEYINPUT1), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT86), .B(new_n289_), .C1(new_n290_), .C2(KEYINPUT1), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n289_), .A2(new_n298_), .A3(KEYINPUT1), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n289_), .B2(KEYINPUT1), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n284_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n303_), .A2(new_n304_), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT88), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n293_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G211gat), .B(G218gat), .Z(new_n315_));
  INV_X1    g114(.A(G197gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT89), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G197gat), .ZN(new_n319_));
  INV_X1    g118(.A(G204gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(G197gat), .B2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n315_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n320_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n326_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(new_n322_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n324_), .A2(new_n327_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n314_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n314_), .A2(new_n333_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n283_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n314_), .A2(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n314_), .A2(new_n333_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n282_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G8gat), .B(G36gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n331_), .B1(new_n226_), .B2(new_n243_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n239_), .B1(new_n241_), .B2(new_n238_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n237_), .B1(new_n221_), .B2(new_n225_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n230_), .A2(new_n210_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n352_), .B1(new_n358_), .B2(new_n331_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n240_), .A2(new_n238_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT78), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n361_), .B(new_n220_), .C1(new_n224_), .C2(new_n223_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n362_), .A2(new_n213_), .B1(new_n242_), .B2(new_n235_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT90), .B1(new_n363_), .B2(new_n331_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n350_), .A2(new_n359_), .A3(new_n364_), .A4(KEYINPUT91), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n358_), .A2(new_n331_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n244_), .B2(new_n332_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n352_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n350_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT91), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n346_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n346_), .A3(new_n368_), .A4(new_n365_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n263_), .A2(new_n266_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n301_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n308_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n292_), .B(new_n377_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n380_), .B(KEYINPUT4), .C1(new_n310_), .C2(new_n267_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n267_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n292_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n380_), .B(new_n382_), .C1(new_n310_), .C2(new_n267_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT33), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n388_), .A2(new_n397_), .A3(new_n389_), .A4(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n381_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n380_), .B(new_n383_), .C1(new_n310_), .C2(new_n267_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n393_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n400_), .B2(new_n393_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n396_), .A2(new_n398_), .B1(new_n404_), .B2(KEYINPUT94), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n399_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n376_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n409_));
  INV_X1    g208(.A(new_n352_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n350_), .A2(new_n364_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n332_), .B1(new_n358_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n412_), .B2(new_n358_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n410_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n366_), .A2(new_n367_), .A3(new_n352_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n388_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n394_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n369_), .A2(new_n372_), .ZN(new_n420_));
  OAI221_X1 g219(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .C1(new_n409_), .C2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n340_), .B1(new_n408_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n374_), .A2(KEYINPUT97), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n369_), .A2(new_n424_), .A3(new_n346_), .A4(new_n372_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n345_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .A4(KEYINPUT27), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT96), .B1(new_n418_), .B2(new_n419_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n388_), .A2(new_n389_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n393_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT96), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n395_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  AND4_X1   g234(.A1(new_n340_), .A2(new_n427_), .A3(new_n429_), .A4(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n277_), .B1(new_n422_), .B2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n427_), .A2(new_n429_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n340_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n269_), .A2(new_n270_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n435_), .A4(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G113gat), .B(G141gat), .Z(new_n442_));
  XOR2_X1   g241(.A(G169gat), .B(G197gat), .Z(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  INV_X1    g243(.A(KEYINPUT73), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT15), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n449_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n447_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n448_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G43gat), .B(G50gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n448_), .A2(new_n449_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT15), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G1gat), .A2(G8gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT14), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n459_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n458_), .A2(new_n459_), .A3(new_n464_), .A4(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n452_), .A2(new_n457_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n455_), .A2(new_n456_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n456_), .A3(new_n455_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n474_), .B2(new_n471_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n446_), .B(KEYINPUT74), .C1(new_n473_), .C2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n472_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n468_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(new_n470_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n469_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n482_), .A3(new_n444_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n482_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT74), .B1(new_n485_), .B2(new_n446_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT75), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n477_), .A2(new_n478_), .B1(new_n481_), .B2(new_n469_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n446_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT75), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n483_), .A4(new_n476_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n437_), .A2(new_n441_), .B1(new_n487_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G230gat), .A2(G233gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT64), .Z(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  AND2_X1   g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT65), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(G85gat), .B2(G92gat), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT10), .B(G99gat), .Z(new_n512_));
  INV_X1    g311(.A(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT66), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n518_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n514_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n497_), .B1(new_n511_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n501_), .A2(new_n506_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n508_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT66), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n528_), .A2(new_n529_), .B1(new_n513_), .B2(new_n512_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n530_), .A3(KEYINPUT67), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT68), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n516_), .A2(new_n518_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537_));
  INV_X1    g336(.A(G99gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n513_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n499_), .A2(new_n500_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT8), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n519_), .A2(new_n520_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n532_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n522_), .A2(new_n531_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n496_), .B1(new_n551_), .B2(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n549_), .A2(KEYINPUT68), .B1(new_n516_), .B2(new_n518_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n546_), .B1(new_n562_), .B2(new_n541_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT8), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n550_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n511_), .A2(new_n521_), .A3(new_n497_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT67), .B1(new_n527_), .B2(new_n530_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n558_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n561_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n559_), .B1(new_n560_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n551_), .A2(new_n558_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n565_), .B(new_n558_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n496_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G120gat), .B(G148gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT70), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n571_), .A2(new_n575_), .A3(new_n583_), .A4(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n571_), .A2(new_n575_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT71), .A3(new_n592_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT34), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT35), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n452_), .A2(new_n457_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n568_), .A2(new_n604_), .B1(new_n601_), .B2(new_n600_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n551_), .A2(new_n470_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT36), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n611_), .B(KEYINPUT36), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT37), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n613_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n619_), .B2(new_n607_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n558_), .A2(new_n480_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n556_), .A2(new_n468_), .A3(new_n557_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(G231gat), .A3(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G127gat), .B(G155gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT17), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n638_), .A3(new_n626_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n628_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n635_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT17), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n633_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n636_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n628_), .B2(new_n639_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n624_), .A2(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n494_), .A2(new_n597_), .A3(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT98), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT98), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n435_), .A2(G1gat), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n650_), .A2(KEYINPUT38), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n437_), .A2(new_n441_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n588_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT13), .B1(new_n585_), .B2(new_n588_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n484_), .A2(new_n486_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n647_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n614_), .A2(new_n617_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n435_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n462_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n657_), .B1(new_n658_), .B2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n655_), .B1(new_n656_), .B2(new_n673_), .ZN(G1324gat));
  INV_X1    g473(.A(new_n438_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n650_), .A2(new_n463_), .A3(new_n675_), .A4(new_n651_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G8gat), .B1(new_n669_), .B2(new_n438_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT100), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(G8gat), .C1(new_n669_), .C2(new_n438_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n679_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n676_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n676_), .B(KEYINPUT40), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(new_n649_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(G15gat), .A3(new_n277_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT101), .ZN(new_n691_));
  OAI21_X1  g490(.A(G15gat), .B1(new_n669_), .B2(new_n277_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT41), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(KEYINPUT41), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n693_), .A3(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n669_), .B2(new_n439_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n439_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n689_), .B2(new_n698_), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n487_), .A2(new_n493_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n667_), .A2(new_n647_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n593_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n659_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n671_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n624_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n624_), .B(KEYINPUT103), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n271_), .A2(new_n276_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n376_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n396_), .A2(new_n398_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n404_), .A2(KEYINPUT94), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n407_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n421_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n439_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n340_), .A2(new_n427_), .A3(new_n429_), .A4(new_n435_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n711_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n441_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n710_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n709_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n665_), .A2(new_n646_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n706_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n722_), .B1(new_n659_), .B2(new_n710_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n725_), .C1(new_n728_), .C2(new_n709_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n671_), .A2(G29gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n705_), .B1(new_n730_), .B2(new_n731_), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n727_), .A2(new_n675_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G36gat), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n438_), .A2(G36gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT104), .B1(new_n703_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n494_), .A2(new_n738_), .A3(new_n702_), .A4(new_n735_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n737_), .A2(KEYINPUT45), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT45), .B1(new_n737_), .B2(new_n739_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n734_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n734_), .A2(KEYINPUT46), .A3(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1329gat));
  NAND4_X1  g546(.A1(new_n727_), .A2(G43gat), .A3(new_n440_), .A4(new_n729_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G43gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n703_), .B2(new_n277_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT106), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n704_), .B2(new_n340_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n340_), .A2(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n730_), .B2(new_n755_), .ZN(G1331gat));
  NAND3_X1  g555(.A1(new_n487_), .A2(new_n646_), .A3(new_n493_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n659_), .A3(new_n668_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n758_), .A2(new_n659_), .A3(KEYINPUT108), .A4(new_n668_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G57gat), .B1(new_n763_), .B2(new_n435_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n648_), .A2(new_n593_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT107), .Z(new_n766_));
  AOI21_X1  g565(.A(new_n664_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n435_), .A2(G57gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT109), .ZN(G1332gat));
  OR3_X1    g570(.A1(new_n768_), .A2(G64gat), .A3(new_n438_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G64gat), .B1(new_n763_), .B2(new_n438_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(KEYINPUT48), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(KEYINPUT48), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(G1333gat));
  OR3_X1    g575(.A1(new_n768_), .A2(G71gat), .A3(new_n277_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n711_), .A3(new_n762_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G71gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT110), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1334gat));
  OR3_X1    g585(.A1(new_n768_), .A2(G78gat), .A3(new_n439_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(new_n340_), .A3(new_n762_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(G78gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(G78gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(G1335gat));
  INV_X1    g591(.A(new_n597_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n767_), .A2(new_n793_), .A3(new_n667_), .A4(new_n647_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n502_), .A3(new_n671_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n662_), .A2(new_n664_), .A3(new_n646_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n724_), .A2(new_n435_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n799_), .B2(new_n502_), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n503_), .A3(new_n675_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n724_), .A2(new_n438_), .A3(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n503_), .ZN(G1337gat));
  NOR2_X1   g602(.A1(new_n724_), .A2(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n711_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n440_), .A2(new_n512_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n805_), .A2(G99gat), .B1(new_n795_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n795_), .A2(new_n513_), .A3(new_n340_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n340_), .B(new_n797_), .C1(new_n728_), .C2(new_n709_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  AND4_X1   g615(.A1(new_n439_), .A2(new_n438_), .A3(new_n671_), .A4(new_n440_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n818_));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n757_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n487_), .A2(new_n493_), .A3(new_n646_), .A4(KEYINPUT111), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n623_), .B2(new_n618_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT112), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT54), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n662_), .A2(new_n829_), .A3(new_n824_), .A4(new_n823_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n496_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n573_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT12), .B1(new_n551_), .B2(new_n558_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n568_), .A2(new_n561_), .A3(new_n569_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n837_));
  AOI21_X1  g636(.A(new_n574_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n836_), .A2(new_n837_), .B1(new_n838_), .B2(new_n832_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n836_), .A2(KEYINPUT55), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n587_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n587_), .B(new_n842_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n663_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n444_), .B1(new_n477_), .B2(new_n472_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n469_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n483_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n589_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n667_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n618_), .A2(new_n623_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n587_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n851_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(KEYINPUT58), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n855_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n862_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n856_), .A2(new_n859_), .A3(new_n864_), .A4(new_n858_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(KEYINPUT57), .A2(new_n854_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n854_), .A2(KEYINPUT57), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n646_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n831_), .B1(new_n868_), .B2(KEYINPUT118), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n847_), .A2(new_n853_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT57), .A3(new_n668_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n860_), .A2(new_n862_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n624_), .A3(new_n865_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n854_), .A2(KEYINPUT57), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n647_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n817_), .B(new_n818_), .C1(new_n869_), .C2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n875_), .A2(KEYINPUT115), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n880_), .A2(new_n866_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n831_), .B1(new_n883_), .B2(new_n646_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(new_n817_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n700_), .B(new_n879_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G113gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n817_), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n889_), .A2(G113gat), .A3(new_n663_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1340gat));
  OAI211_X1 g690(.A(new_n793_), .B(new_n879_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G120gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n662_), .A2(KEYINPUT60), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n894_), .B(KEYINPUT60), .S(G120gat), .Z(new_n895_));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1341gat));
  OAI211_X1 g696(.A(new_n646_), .B(new_n879_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G127gat), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n889_), .A2(G127gat), .A3(new_n647_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  OAI211_X1 g700(.A(new_n624_), .B(new_n879_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G134gat), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n889_), .A2(G134gat), .A3(new_n668_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1343gat));
  NAND4_X1  g704(.A1(new_n277_), .A2(new_n438_), .A3(new_n340_), .A4(new_n671_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT119), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n884_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n663_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT120), .B(G141gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n908_), .A2(new_n597_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT121), .B(G148gat), .Z(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1345gat));
  NOR2_X1   g713(.A1(new_n908_), .A2(new_n647_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT61), .B(G155gat), .Z(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  INV_X1    g716(.A(new_n908_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n918_), .A2(G162gat), .A3(new_n710_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G162gat), .B1(new_n918_), .B2(new_n667_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1347gat));
  NOR3_X1   g720(.A1(new_n277_), .A2(new_n438_), .A3(new_n671_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n439_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n826_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n868_), .A2(KEYINPUT118), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n663_), .B(new_n925_), .C1(new_n927_), .C2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT123), .B1(new_n929_), .B2(new_n207_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n925_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n664_), .B(new_n931_), .C1(new_n869_), .C2(new_n878_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n932_), .A2(new_n933_), .A3(G169gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(KEYINPUT62), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n233_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n932_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n932_), .B2(G169gat), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n935_), .A2(new_n940_), .ZN(G1348gat));
  AOI21_X1  g740(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n942_));
  AOI21_X1  g741(.A(G176gat), .B1(new_n942_), .B2(new_n593_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n884_), .A2(new_n439_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n924_), .A2(G176gat), .A3(new_n793_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n943_), .A2(new_n946_), .ZN(G1349gat));
  AND4_X1   g746(.A1(new_n439_), .A2(new_n884_), .A3(new_n646_), .A4(new_n924_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(G183gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n647_), .A2(new_n204_), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n942_), .A2(KEYINPUT124), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(KEYINPUT124), .B1(new_n942_), .B2(new_n950_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n949_), .A2(new_n951_), .A3(new_n952_), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n942_), .A2(new_n205_), .A3(new_n667_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n942_), .A2(new_n624_), .ZN(new_n955_));
  INV_X1    g754(.A(G190gat), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G1351gat));
  NOR4_X1   g756(.A1(new_n711_), .A2(new_n438_), .A3(new_n439_), .A4(new_n671_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n884_), .A2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n316_), .A2(KEYINPUT125), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n316_), .A2(KEYINPUT125), .ZN(new_n962_));
  AOI22_X1  g761(.A1(new_n960_), .A2(new_n664_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n959_), .A2(new_n663_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n962_), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n959_), .A2(new_n597_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n320_), .ZN(G1353gat));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n959_), .A2(new_n647_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n968_), .B1(new_n969_), .B2(new_n971_), .ZN(new_n972_));
  OAI211_X1 g771(.A(KEYINPUT126), .B(new_n970_), .C1(new_n959_), .C2(new_n647_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT63), .B(G211gat), .Z(new_n974_));
  AOI22_X1  g773(.A1(new_n972_), .A2(new_n973_), .B1(new_n969_), .B2(new_n974_), .ZN(G1354gat));
  OR3_X1    g774(.A1(new_n959_), .A2(G218gat), .A3(new_n668_), .ZN(new_n976_));
  OAI21_X1  g775(.A(G218gat), .B1(new_n959_), .B2(new_n855_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1355gat));
endmodule


