//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT105), .B(KEYINPUT20), .Z(new_n206_));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT91), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT89), .B(G197gat), .Z(new_n215_));
  INV_X1    g014(.A(G204gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n212_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(G204gat), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n216_), .B2(G197gat), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT21), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n216_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n218_), .B1(new_n229_), .B2(new_n213_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n212_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n212_), .A2(KEYINPUT92), .A3(new_n228_), .A4(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n219_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT26), .B(G190gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT96), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT25), .B(G183gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT23), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n242_), .B1(new_n246_), .B2(KEYINPUT81), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT24), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n246_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT80), .B(G176gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n257_), .A2(new_n258_), .B1(G169gat), .B2(G176gat), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n240_), .A2(new_n255_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n206_), .B1(new_n235_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n219_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n217_), .A2(new_n218_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT92), .B1(new_n263_), .B2(new_n228_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n234_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n254_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n239_), .A2(new_n236_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI221_X1 g068(.A(new_n242_), .B1(G183gat), .B2(G190gat), .C1(new_n246_), .C2(KEYINPUT81), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n248_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT22), .B1(new_n248_), .B2(KEYINPUT79), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n257_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n252_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n269_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n266_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n205_), .B1(new_n261_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT97), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n240_), .A2(new_n255_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n259_), .A2(new_n256_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n266_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT97), .B1(new_n235_), .B2(new_n260_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n285_));
  INV_X1    g084(.A(new_n276_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n235_), .B2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n283_), .A2(new_n284_), .A3(new_n287_), .A4(new_n205_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT106), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n278_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n284_), .A2(new_n287_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT106), .A3(new_n205_), .A4(new_n283_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT100), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G8gat), .B(G36gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT99), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n297_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT108), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(KEYINPUT108), .A3(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n283_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n204_), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n285_), .B(new_n204_), .C1(new_n235_), .C2(new_n260_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n277_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n300_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n306_), .A2(new_n204_), .B1(new_n277_), .B2(new_n308_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT101), .B1(new_n314_), .B2(new_n310_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n311_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n314_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n317_), .A2(KEYINPUT101), .A3(new_n300_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n305_), .A2(new_n313_), .B1(new_n319_), .B2(new_n312_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT0), .ZN(new_n322_));
  INV_X1    g121(.A(G57gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n330_), .A2(KEYINPUT83), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(KEYINPUT83), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n334_));
  INV_X1    g133(.A(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n339_), .A2(KEYINPUT86), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT87), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT86), .B1(new_n339_), .B2(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(KEYINPUT85), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n340_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n342_), .A2(KEYINPUT87), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n338_), .B1(new_n346_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n339_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n351_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n333_), .A2(new_n336_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n337_), .B(KEYINPUT1), .Z(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n328_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n359_), .B(new_n337_), .C1(new_n345_), .C2(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n351_), .A3(new_n357_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(KEYINPUT88), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G127gat), .B(G134gat), .Z(new_n367_));
  XOR2_X1   g166(.A(G113gat), .B(G120gat), .Z(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n369_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n365_), .A3(new_n363_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n372_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n327_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT107), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n370_), .A2(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT4), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n370_), .A2(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n378_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n326_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT107), .B(new_n327_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT28), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n362_), .A2(new_n366_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n392_), .ZN(new_n396_));
  AOI211_X1 g195(.A(KEYINPUT29), .B(new_n396_), .C1(new_n362_), .C2(new_n366_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n394_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n399_));
  OAI211_X1 g198(.A(G228gat), .B(G233gat), .C1(new_n235_), .C2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n362_), .A2(KEYINPUT29), .A3(new_n366_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n266_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n400_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n398_), .B1(new_n406_), .B2(KEYINPUT94), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n266_), .B(new_n402_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n400_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n400_), .B(new_n408_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n410_), .A2(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n409_), .A2(KEYINPUT95), .A3(new_n408_), .A4(new_n400_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(KEYINPUT93), .A3(new_n412_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n404_), .A2(new_n418_), .A3(new_n405_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n398_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n269_), .B(KEYINPUT30), .C1(new_n271_), .C2(new_n275_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n274_), .A2(new_n252_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n270_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT30), .B1(new_n431_), .B2(new_n269_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n276_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n427_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n428_), .A3(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n433_), .A2(new_n373_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n373_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n424_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n369_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n373_), .A3(new_n437_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n423_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n444_), .A3(KEYINPUT82), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n421_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n416_), .A2(new_n445_), .A3(new_n420_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n390_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n300_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT104), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n293_), .A2(new_n454_), .B1(new_n455_), .B2(new_n314_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n389_), .A3(new_n388_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n326_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT33), .B1(new_n458_), .B2(KEYINPUT102), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT102), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n372_), .A2(new_n375_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n379_), .B1(new_n462_), .B2(new_n378_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n460_), .B(new_n461_), .C1(new_n463_), .C2(new_n326_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n382_), .A2(new_n376_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n327_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n383_), .A2(new_n384_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT103), .B1(new_n467_), .B2(new_n376_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT103), .B(new_n376_), .C1(new_n372_), .C2(new_n375_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n459_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n457_), .B1(new_n319_), .B2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n440_), .A2(new_n444_), .A3(KEYINPUT82), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT82), .B1(new_n440_), .B2(new_n444_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n421_), .A2(new_n476_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n320_), .A2(new_n452_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  INV_X1    g279(.A(G43gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G36gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G29gat), .ZN(new_n484_));
  INV_X1    g283(.A(G29gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G36gat), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(new_n486_), .A3(new_n481_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n482_), .A2(new_n487_), .A3(KEYINPUT72), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G43gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n481_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G50gat), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n488_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT72), .B1(new_n482_), .B2(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n489_), .ZN(new_n497_));
  AOI21_X1  g296(.A(G50gat), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n479_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(G50gat), .A3(new_n497_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT15), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G1gat), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT74), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(KEYINPUT14), .C1(new_n504_), .C2(new_n505_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G1gat), .B(G8gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n500_), .A2(new_n501_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n495_), .A2(new_n498_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n513_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n519_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G169gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n225_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT78), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n527_), .B(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n478_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT77), .ZN(new_n537_));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  XNOR2_X1  g338(.A(G183gat), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT75), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n513_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n545_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT11), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n545_), .B(new_n546_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n555_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n543_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n541_), .B(new_n542_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n557_), .A2(new_n559_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G85gat), .B(G92gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT6), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n568_));
  NOR3_X1   g367(.A1(KEYINPUT64), .A2(G99gat), .A3(G106gat), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n567_), .B(new_n568_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  NOR4_X1   g370(.A1(KEYINPUT64), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT65), .B(new_n564_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT66), .B(new_n564_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(KEYINPUT8), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT10), .B(G99gat), .Z(new_n578_));
  INV_X1    g377(.A(G106gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n564_), .A2(KEYINPUT9), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n567_), .A2(new_n568_), .ZN(new_n582_));
  INV_X1    g381(.A(G92gat), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n325_), .A2(new_n583_), .A3(KEYINPUT9), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT8), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n574_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n577_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n503_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n593_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n587_), .A2(new_n585_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n522_), .A2(new_n597_), .A3(new_n577_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n589_), .A2(new_n595_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n588_), .B2(new_n516_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n499_), .A2(new_n502_), .B1(new_n597_), .B2(new_n577_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n594_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT36), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n602_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(KEYINPUT73), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n608_), .B(new_n610_), .C1(KEYINPUT73), .C2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n563_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT68), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n555_), .B1(new_n597_), .B2(new_n577_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n575_), .A2(KEYINPUT8), .A3(new_n576_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n587_), .A2(new_n585_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n556_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n619_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT68), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(KEYINPUT12), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n577_), .A2(new_n585_), .A3(new_n555_), .A4(new_n587_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n620_), .A2(new_n625_), .A3(new_n626_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n627_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT70), .ZN(new_n635_));
  XOR2_X1   g434(.A(G176gat), .B(G204gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  NAND3_X1  g438(.A1(new_n630_), .A2(new_n633_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT71), .ZN(new_n643_));
  OAI22_X1  g442(.A1(new_n641_), .A2(new_n642_), .B1(new_n643_), .B2(KEYINPUT13), .ZN(new_n644_));
  INV_X1    g443(.A(new_n642_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n640_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n616_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n535_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n390_), .A2(new_n504_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n202_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT111), .Z(new_n653_));
  INV_X1    g452(.A(new_n611_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n648_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n534_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n478_), .A2(new_n654_), .A3(new_n657_), .A4(new_n563_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n504_), .B1(new_n658_), .B2(new_n390_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT110), .Z(new_n660_));
  NOR3_X1   g459(.A1(new_n650_), .A2(new_n202_), .A3(new_n651_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n653_), .A2(new_n660_), .A3(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n320_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n505_), .B1(new_n658_), .B2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT112), .B(KEYINPUT39), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n650_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n505_), .A3(new_n665_), .ZN(new_n670_));
  OR2_X1    g469(.A1(KEYINPUT112), .A2(KEYINPUT39), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n668_), .B(new_n670_), .C1(new_n666_), .C2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n666_), .A2(new_n671_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT40), .A3(new_n668_), .A4(new_n670_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n658_), .B2(new_n476_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n669_), .A2(new_n678_), .A3(new_n476_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n680_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n658_), .B2(new_n421_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT42), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n669_), .A2(new_n685_), .A3(new_n421_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n563_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n655_), .A2(new_n611_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n535_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n388_), .A2(new_n389_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n485_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n657_), .A2(new_n690_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n473_), .A2(new_n477_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n412_), .A2(new_n413_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n404_), .A2(new_n411_), .A3(new_n405_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n415_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n419_), .A2(new_n398_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n700_), .A2(new_n407_), .B1(new_n701_), .B2(new_n417_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n451_), .B1(new_n702_), .B2(new_n476_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n293_), .B2(new_n300_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n302_), .B(new_n310_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n313_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n315_), .A2(new_n311_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n315_), .A2(new_n311_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n312_), .A3(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n703_), .A2(new_n706_), .A3(new_n693_), .A4(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n697_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n613_), .A2(new_n615_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n696_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n697_), .B2(new_n710_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT44), .B(new_n695_), .C1(new_n714_), .C2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(G29gat), .A3(new_n390_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n695_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n613_), .A2(new_n615_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT114), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n478_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n717_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT44), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n694_), .B1(new_n719_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT115), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n694_), .C1(new_n719_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1328gat));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n320_), .B1(new_n725_), .B2(KEYINPUT44), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n714_), .A2(new_n717_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n720_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n483_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n665_), .A2(new_n483_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT45), .B1(new_n692_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n740_));
  INV_X1    g539(.A(new_n738_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n535_), .A2(new_n740_), .A3(new_n691_), .A4(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n732_), .B1(new_n737_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n718_), .A2(new_n665_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G36gat), .B1(new_n726_), .B2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(KEYINPUT46), .A3(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1329gat));
  OAI21_X1  g548(.A(new_n481_), .B1(new_n692_), .B2(new_n449_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n481_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n718_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n726_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g553(.A(new_n692_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G50gat), .B1(new_n755_), .B2(new_n421_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n718_), .A2(G50gat), .A3(new_n421_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n736_), .ZN(G1331gat));
  XNOR2_X1  g557(.A(new_n527_), .B(new_n532_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n655_), .A2(new_n690_), .ZN(new_n760_));
  OR4_X1    g559(.A1(new_n478_), .A2(new_n654_), .A3(new_n759_), .A4(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n693_), .ZN(new_n762_));
  NOR4_X1   g561(.A1(new_n478_), .A2(new_n759_), .A3(new_n721_), .A4(new_n760_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n323_), .A3(new_n390_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n766_), .A3(new_n665_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G64gat), .B1(new_n761_), .B2(new_n320_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n772_), .A3(new_n476_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n761_), .B2(new_n449_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n763_), .A2(new_n778_), .A3(new_n421_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G78gat), .B1(new_n761_), .B2(new_n702_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(G78gat), .C1(new_n761_), .C2(new_n702_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n781_), .A2(KEYINPUT50), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT50), .B1(new_n781_), .B2(new_n783_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n779_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n478_), .A2(new_n759_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n690_), .A2(new_n648_), .A3(new_n611_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n325_), .A3(new_n390_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n723_), .A2(new_n724_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n690_), .A2(new_n648_), .A3(new_n759_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(new_n390_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(new_n325_), .ZN(G1336gat));
  NAND3_X1  g595(.A1(new_n790_), .A2(new_n583_), .A3(new_n665_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n794_), .A2(new_n665_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n583_), .ZN(G1337gat));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n445_), .A2(new_n578_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n789_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n792_), .A2(new_n476_), .A3(new_n793_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(G99gat), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n790_), .A2(new_n579_), .A3(new_n421_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n421_), .B(new_n793_), .C1(new_n714_), .C2(new_n717_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G106gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G106gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT53), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n808_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n320_), .A2(new_n390_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n451_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n525_), .A2(new_n518_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n531_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n518_), .B(new_n517_), .C1(new_n503_), .C2(new_n514_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n515_), .A2(new_n523_), .A3(new_n519_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT120), .A3(new_n531_), .A4(new_n822_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n825_), .A2(new_n827_), .B1(new_n530_), .B2(new_n527_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n640_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n623_), .A2(new_n624_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n830_), .A2(new_n617_), .B1(KEYINPUT12), .B2(new_n618_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n625_), .A4(new_n629_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n620_), .A2(new_n625_), .A3(new_n627_), .A4(new_n626_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n632_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n835_));
  NAND2_X1  g634(.A1(new_n630_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n639_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(KEYINPUT56), .A3(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n829_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n721_), .B1(new_n843_), .B2(KEYINPUT58), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n828_), .A2(new_n640_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n837_), .A2(KEYINPUT56), .A3(new_n838_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n838_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n845_), .B(KEYINPUT58), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n534_), .A2(new_n641_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n645_), .A2(new_n640_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n828_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n654_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n844_), .A2(new_n849_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n759_), .A2(new_n640_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n853_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n611_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n563_), .B1(new_n855_), .B2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n712_), .A2(new_n690_), .A3(new_n648_), .A4(new_n534_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT118), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n616_), .A2(new_n865_), .A3(new_n534_), .A4(new_n648_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n864_), .A2(KEYINPUT54), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n864_), .B2(new_n866_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n820_), .B1(new_n862_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870_), .B2(new_n759_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n712_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n860_), .A2(new_n859_), .B1(new_n875_), .B2(new_n848_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n854_), .A2(KEYINPUT57), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n690_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n864_), .A2(new_n866_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n864_), .A2(KEYINPUT54), .A3(new_n866_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n872_), .B(new_n819_), .C1(new_n878_), .C2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n819_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n759_), .A2(KEYINPUT122), .A3(G113gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(KEYINPUT122), .B2(G113gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n871_), .B1(new_n890_), .B2(new_n892_), .ZN(G1340gat));
  INV_X1    g692(.A(G120gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n648_), .B2(KEYINPUT60), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n870_), .B(new_n895_), .C1(KEYINPUT60), .C2(new_n894_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n884_), .A2(new_n655_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n894_), .ZN(G1341gat));
  AOI21_X1  g698(.A(G127gat), .B1(new_n870_), .B2(new_n690_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n690_), .A2(G127gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT123), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n890_), .B2(new_n902_), .ZN(G1342gat));
  AOI21_X1  g702(.A(G134gat), .B1(new_n870_), .B2(new_n654_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT124), .B(G134gat), .Z(new_n905_));
  NOR2_X1   g704(.A1(new_n712_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n890_), .B2(new_n906_), .ZN(G1343gat));
  AOI211_X1 g706(.A(new_n450_), .B(new_n818_), .C1(new_n862_), .C2(new_n869_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n759_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n655_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n690_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n913_), .B(new_n915_), .ZN(G1346gat));
  AOI21_X1  g715(.A(G162gat), .B1(new_n908_), .B2(new_n654_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n713_), .A2(G162gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n908_), .B2(new_n918_), .ZN(G1347gat));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n862_), .A2(new_n869_), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n320_), .A2(new_n390_), .A3(new_n449_), .A4(new_n421_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n534_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n920_), .B1(new_n924_), .B2(new_n248_), .ZN(new_n925_));
  OAI211_X1 g724(.A(KEYINPUT62), .B(G169gat), .C1(new_n923_), .C2(new_n534_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n258_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(G1348gat));
  NOR3_X1   g727(.A1(new_n923_), .A2(new_n249_), .A3(new_n648_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n923_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n655_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n257_), .B2(new_n931_), .ZN(G1349gat));
  AOI21_X1  g731(.A(G183gat), .B1(new_n930_), .B2(new_n690_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n923_), .A2(new_n239_), .A3(new_n563_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n923_), .B2(new_n712_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n654_), .A2(new_n238_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n923_), .B2(new_n937_), .ZN(G1351gat));
  INV_X1    g737(.A(new_n450_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n320_), .A2(new_n390_), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n921_), .A2(new_n939_), .A3(new_n759_), .A4(new_n940_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n941_), .A2(KEYINPUT126), .A3(new_n225_), .ZN(new_n942_));
  AOI21_X1  g741(.A(KEYINPUT126), .B1(new_n941_), .B2(new_n225_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n225_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n942_), .A2(new_n943_), .A3(new_n944_), .ZN(G1352gat));
  NAND3_X1  g744(.A1(new_n921_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n648_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n216_), .ZN(G1353gat));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949_));
  INV_X1    g748(.A(G211gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n690_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n946_), .A2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n950_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT127), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n952_), .B(new_n954_), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n946_), .B2(new_n712_), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n611_), .A2(G218gat), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n946_), .B2(new_n957_), .ZN(G1355gat));
endmodule


