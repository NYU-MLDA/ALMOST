//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G50gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT74), .ZN(new_n209_));
  INV_X1    g008(.A(G15gat), .ZN(new_n210_));
  INV_X1    g009(.A(G22gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G15gat), .A2(G22gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G1gat), .A2(G8gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n212_), .A2(new_n213_), .B1(KEYINPUT14), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n209_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G229gat), .A2(G233gat), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n205_), .A2(new_n216_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n205_), .B(new_n216_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G229gat), .A3(G233gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G113gat), .B(G141gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G197gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n222_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(KEYINPUT75), .A3(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G8gat), .B(G36gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G64gat), .B(G92gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G211gat), .B(G218gat), .Z(new_n242_));
  INV_X1    g041(.A(G204gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(KEYINPUT85), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT85), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n226_), .A2(G204gat), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT21), .B(new_n242_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT86), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G197gat), .A2(G204gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT85), .B(G197gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT21), .B(new_n251_), .C1(new_n252_), .C2(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  INV_X1    g053(.A(new_n248_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n255_), .C1(new_n252_), .C2(new_n243_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n242_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n255_), .B1(new_n252_), .B2(new_n243_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT21), .A4(new_n242_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n250_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT76), .B(G183gat), .ZN(new_n263_));
  INV_X1    g062(.A(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT23), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT81), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n266_), .B2(KEYINPUT23), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n265_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT78), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G169gat), .A3(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT22), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(G169gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n279_), .B(new_n282_), .C1(new_n283_), .C2(new_n280_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n273_), .A2(new_n278_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n293_), .B2(KEYINPUT25), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT77), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G190gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(KEYINPUT77), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n289_), .B(KEYINPUT79), .C1(new_n294_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n267_), .A2(new_n269_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n295_), .B2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n308_), .B2(new_n305_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n290_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n263_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n288_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n304_), .B1(new_n313_), .B2(KEYINPUT79), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n262_), .B(new_n286_), .C1(new_n302_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT87), .Z(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT19), .Z(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  INV_X1    g118(.A(new_n272_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n301_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT81), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n296_), .A2(new_n307_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n296_), .B2(new_n307_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n323_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n287_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n303_), .B1(new_n328_), .B2(new_n274_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n283_), .A2(new_n279_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n278_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n250_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n319_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n315_), .A2(new_n318_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n286_), .B1(new_n314_), .B2(new_n302_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n241_), .B(new_n337_), .C1(new_n340_), .C2(new_n318_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n241_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n335_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n338_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n318_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n315_), .A2(new_n318_), .A3(new_n336_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n318_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n289_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n303_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n321_), .B1(new_n313_), .B2(KEYINPUT79), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n262_), .B1(new_n355_), .B2(new_n286_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n356_), .B2(new_n338_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n357_), .A2(KEYINPUT90), .A3(new_n241_), .A4(new_n337_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n343_), .A2(new_n349_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  AND2_X1   g159(.A1(G127gat), .A2(G134gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(G113gat), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G127gat), .ZN(new_n364_));
  INV_X1    g163(.A(G134gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G113gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G127gat), .A2(G134gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n363_), .A2(new_n369_), .A3(G120gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(G120gat), .B1(new_n363_), .B2(new_n369_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373_));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT83), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n374_), .B2(KEYINPUT1), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381_));
  INV_X1    g180(.A(G141gat), .ZN(new_n382_));
  INV_X1    g181(.A(G148gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n384_), .A2(new_n387_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n376_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n390_), .A2(new_n391_), .B1(new_n373_), .B2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n372_), .B(new_n380_), .C1(new_n375_), .C2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n363_), .A2(new_n369_), .ZN(new_n395_));
  INV_X1    g194(.A(G120gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n363_), .A2(new_n369_), .A3(G120gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n373_), .A2(new_n392_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n375_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n380_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n394_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n394_), .A2(new_n404_), .A3(KEYINPUT92), .A4(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n394_), .A2(new_n404_), .A3(KEYINPUT4), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n400_), .A2(new_n401_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n374_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n380_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n399_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n405_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n415_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n410_), .A2(new_n415_), .A3(new_n423_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n416_), .A2(new_n421_), .A3(new_n405_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n415_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n394_), .A2(new_n404_), .A3(new_n422_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n359_), .A2(new_n360_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G78gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n335_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n418_), .A2(new_n443_), .A3(new_n444_), .A4(new_n380_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n380_), .C1(new_n393_), .C2(new_n375_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT28), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n419_), .A2(KEYINPUT29), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n335_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n440_), .A2(new_n445_), .A3(new_n447_), .A4(new_n441_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n438_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n452_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n451_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n437_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n318_), .B1(new_n356_), .B2(new_n338_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n315_), .A2(new_n350_), .A3(new_n336_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n410_), .A2(new_n423_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n428_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n469_), .B2(new_n426_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n461_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n343_), .A2(new_n349_), .A3(new_n358_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n431_), .A2(new_n426_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n424_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT93), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n433_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n339_), .A2(KEYINPUT30), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n355_), .A2(new_n478_), .A3(new_n286_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT82), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G43gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT31), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n478_), .B1(new_n355_), .B2(new_n286_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT30), .B(new_n285_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n491_));
  INV_X1    g290(.A(new_n485_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n486_), .A2(new_n493_), .A3(new_n399_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n399_), .B1(new_n486_), .B2(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT82), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n480_), .A2(KEYINPUT31), .A3(new_n485_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n372_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n486_), .A2(new_n493_), .A3(new_n399_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n476_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n469_), .A2(new_n426_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT27), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n472_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n350_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n315_), .A2(new_n350_), .A3(new_n336_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n241_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n513_), .B2(new_n349_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n344_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT27), .B1(new_n515_), .B2(KEYINPUT94), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n514_), .A2(new_n516_), .A3(KEYINPUT95), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n241_), .B1(new_n357_), .B2(new_n337_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT94), .B1(new_n515_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n508_), .B1(new_n513_), .B2(new_n510_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n507_), .B(new_n509_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n461_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n505_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT95), .B1(new_n514_), .B2(new_n516_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n520_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n526_), .A2(new_n527_), .B1(new_n508_), .B2(new_n472_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n496_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n501_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n506_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n461_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n236_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT96), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT10), .B(G99gat), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n435_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT64), .B(G92gat), .Z(new_n543_));
  INV_X1    g342(.A(KEYINPUT9), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(G85gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G85gat), .B(G92gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(new_n544_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT66), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT66), .ZN(new_n553_));
  NOR2_X1   g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n540_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT8), .ZN(new_n557_));
  INV_X1    g356(.A(new_n547_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT67), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n550_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566_));
  AND3_X1   g365(.A1(new_n565_), .A2(KEYINPUT11), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n565_), .B2(KEYINPUT11), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n565_), .A2(KEYINPUT11), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n570_), .B(new_n550_), .C1(new_n561_), .C2(new_n560_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n537_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT69), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT12), .B1(new_n562_), .B2(new_n571_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n573_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT70), .B1(new_n546_), .B2(new_n548_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n545_), .A2(new_n542_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n586_));
  INV_X1    g385(.A(new_n548_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n540_), .A4(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n560_), .A2(new_n561_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT12), .B(new_n571_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n537_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n575_), .A2(new_n580_), .A3(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n575_), .A2(new_n592_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n580_), .B(KEYINPUT72), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n536_), .B(new_n593_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n575_), .A2(new_n580_), .A3(new_n592_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n596_), .B1(new_n575_), .B2(new_n592_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT13), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G134gat), .ZN(new_n603_));
  INV_X1    g402(.A(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n207_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n562_), .A2(new_n205_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(KEYINPUT35), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n608_), .A2(new_n609_), .A3(new_n614_), .A4(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n607_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(new_n605_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n607_), .A3(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(KEYINPUT73), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(KEYINPUT37), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n619_), .B(new_n620_), .C1(KEYINPUT73), .C2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n570_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n216_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G183gat), .ZN(new_n633_));
  INV_X1    g432(.A(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n629_), .A2(new_n630_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(KEYINPUT17), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n626_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n535_), .A2(new_n601_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT97), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n535_), .A2(new_n644_), .A3(new_n601_), .A4(new_n641_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G1gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n506_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n601_), .A2(new_n235_), .A3(new_n639_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n621_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n507_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n648_), .A2(new_n649_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n650_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(G8gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n528_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n643_), .A2(new_n661_), .A3(new_n662_), .A4(new_n645_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G8gat), .B1(new_n657_), .B2(new_n528_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT99), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(G8gat), .C1(new_n657_), .C2(new_n528_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(KEYINPUT39), .A3(new_n667_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n663_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT100), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n663_), .A2(new_n670_), .A3(new_n674_), .A4(new_n671_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n673_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n673_), .B2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1325gat));
  INV_X1    g477(.A(new_n504_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n646_), .A2(new_n210_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G15gat), .B1(new_n657_), .B2(new_n504_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT41), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1326gat));
  NAND3_X1  g482(.A1(new_n646_), .A2(new_n211_), .A3(new_n461_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G22gat), .B1(new_n657_), .B2(new_n532_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT42), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n621_), .A2(new_n639_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n535_), .A2(new_n601_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n506_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n532_), .B1(new_n528_), .B2(new_n507_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n476_), .A2(new_n504_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n533_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT101), .B(new_n533_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n626_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n626_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT43), .B1(new_n525_), .B2(new_n533_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT102), .A3(new_n626_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n699_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n601_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n236_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n708_), .A4(new_n640_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n709_), .A2(G29gat), .A3(new_n506_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n703_), .A2(new_n705_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(new_n640_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n691_), .B1(new_n710_), .B2(new_n715_), .ZN(G1328gat));
  OR3_X1    g515(.A1(new_n689_), .A2(G36gat), .A3(new_n528_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n709_), .A2(new_n662_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT102), .B1(new_n704_), .B2(new_n626_), .ZN(new_n721_));
  AND4_X1   g520(.A1(KEYINPUT102), .A2(new_n694_), .A3(new_n626_), .A4(new_n700_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n639_), .B1(new_n723_), .B2(new_n699_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n724_), .B2(new_n708_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n719_), .B(G36gat), .C1(new_n720_), .C2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n715_), .A2(new_n662_), .A3(new_n709_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n719_), .B1(new_n728_), .B2(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n718_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n718_), .B(KEYINPUT46), .C1(new_n727_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  OAI21_X1  g533(.A(new_n203_), .B1(new_n689_), .B2(new_n504_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n715_), .A2(G43gat), .A3(new_n679_), .A4(new_n709_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n690_), .B2(new_n461_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n715_), .A2(G50gat), .A3(new_n461_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n709_), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n601_), .A2(new_n235_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n656_), .A2(new_n639_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n506_), .B2(G57gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n694_), .A2(new_n744_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n641_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT105), .Z(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n506_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n752_));
  INV_X1    g551(.A(G57gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(G1332gat));
  OAI21_X1  g553(.A(G64gat), .B1(new_n745_), .B2(new_n528_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT48), .ZN(new_n756_));
  INV_X1    g555(.A(new_n751_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n528_), .A2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n745_), .B2(new_n504_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n504_), .A2(G71gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n757_), .B2(new_n762_), .ZN(G1334gat));
  OAI21_X1  g562(.A(G78gat), .B1(new_n745_), .B2(new_n532_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT50), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n532_), .A2(G78gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n757_), .B2(new_n766_), .ZN(G1335gat));
  OR2_X1    g566(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n601_), .A2(new_n235_), .A3(new_n639_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n507_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n749_), .A2(new_n688_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT107), .Z(new_n774_));
  INV_X1    g573(.A(G85gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n506_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT109), .ZN(G1336gat));
  AOI21_X1  g577(.A(G92gat), .B1(new_n774_), .B2(new_n662_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n771_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n662_), .A2(new_n543_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n771_), .B2(new_n504_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n774_), .A2(new_n541_), .A3(new_n679_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1338gat));
  NAND4_X1  g588(.A1(new_n706_), .A2(new_n640_), .A3(new_n461_), .A4(new_n744_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT111), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n774_), .A2(new_n435_), .A3(new_n461_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(KEYINPUT111), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n795_), .A2(new_n796_), .A3(new_n801_), .A4(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n679_), .A2(new_n506_), .A3(new_n528_), .A4(new_n532_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT116), .Z(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT12), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n556_), .A2(new_n559_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT8), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n549_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n811_), .B2(new_n570_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n591_), .A2(new_n812_), .A3(new_n573_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n537_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n806_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n813_), .A2(new_n814_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n813_), .A2(new_n806_), .A3(new_n814_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n595_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n221_), .A2(new_n218_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n217_), .A2(new_n219_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n227_), .B(new_n821_), .C1(new_n822_), .C2(new_n218_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n230_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n595_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n820_), .A2(new_n593_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT58), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n537_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n592_), .B1(new_n830_), .B2(new_n806_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n818_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n833_), .B2(new_n595_), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT56), .B(new_n596_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT114), .A3(new_n593_), .A4(new_n824_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n626_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT115), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n836_), .A2(KEYINPUT58), .A3(new_n593_), .A4(new_n824_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n842_), .A3(new_n626_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n820_), .A2(new_n235_), .A3(new_n593_), .A4(new_n826_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n824_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n621_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT57), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n639_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n601_), .A2(new_n236_), .A3(new_n639_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT112), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n623_), .A2(new_n625_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n601_), .A2(new_n855_), .A3(new_n236_), .A4(new_n639_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .A4(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT54), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n852_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(KEYINPUT113), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT113), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(KEYINPUT54), .A3(new_n857_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n805_), .B1(new_n850_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n235_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(KEYINPUT59), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n858_), .B(new_n861_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n848_), .B(KEYINPUT57), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n842_), .B1(new_n838_), .B2(new_n626_), .ZN(new_n870_));
  AOI211_X1 g669(.A(KEYINPUT115), .B(new_n854_), .C1(new_n829_), .C2(new_n837_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n872_), .B2(new_n841_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n868_), .B1(new_n873_), .B2(new_n639_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n805_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n867_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n236_), .A2(new_n367_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n866_), .B1(new_n877_), .B2(new_n878_), .ZN(G1340gat));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880_));
  AOI21_X1  g679(.A(G120gat), .B1(new_n707_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n396_), .A2(KEYINPUT60), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n864_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n867_), .A2(new_n876_), .A3(new_n707_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G120gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1341gat));
  NAND2_X1  g687(.A1(new_n639_), .A2(G127gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT118), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n867_), .A2(new_n876_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n364_), .B1(new_n864_), .B2(new_n640_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(KEYINPUT119), .A3(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1342gat));
  OAI21_X1  g696(.A(new_n365_), .B1(new_n864_), .B2(new_n621_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n898_), .A2(KEYINPUT120), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(KEYINPUT120), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n854_), .A2(new_n365_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT121), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n899_), .A2(new_n900_), .B1(new_n877_), .B2(new_n902_), .ZN(G1343gat));
  OAI211_X1 g702(.A(new_n461_), .B(new_n504_), .C1(new_n850_), .C2(new_n863_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n904_), .A2(new_n507_), .A3(new_n662_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n235_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n707_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n639_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  AOI21_X1  g711(.A(G162gat), .B1(new_n905_), .B2(new_n655_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n854_), .A2(new_n604_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(G1347gat));
  NAND3_X1  g714(.A1(new_n662_), .A2(new_n532_), .A3(new_n531_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n235_), .B(new_n917_), .C1(new_n850_), .C2(new_n863_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(KEYINPUT122), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n918_), .A2(new_n921_), .A3(G169gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n850_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n916_), .B1(new_n926_), .B2(new_n868_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(new_n235_), .A3(new_n283_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n920_), .A2(KEYINPUT62), .A3(new_n922_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n925_), .A2(new_n928_), .A3(new_n929_), .ZN(G1348gat));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n707_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n874_), .A2(new_n639_), .A3(new_n917_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT123), .B1(new_n933_), .B2(new_n323_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  INV_X1    g734(.A(new_n323_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n927_), .A2(new_n935_), .A3(new_n639_), .A4(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n933_), .B(KEYINPUT124), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n263_), .B2(new_n939_), .ZN(G1350gat));
  OAI211_X1 g739(.A(new_n927_), .B(new_n655_), .C1(new_n326_), .C2(new_n325_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n927_), .A2(new_n626_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n943_), .B2(new_n264_), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n528_), .A2(new_n506_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n874_), .A2(new_n461_), .A3(new_n504_), .A4(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n236_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n226_), .ZN(G1352gat));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n601_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(new_n243_), .ZN(G1353gat));
  AOI21_X1  g749(.A(new_n679_), .B1(new_n926_), .B2(new_n868_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n951_), .A2(new_n639_), .A3(new_n461_), .A4(new_n945_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT63), .B(G211gat), .Z(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT125), .B1(new_n952_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n946_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n956_), .A2(new_n957_), .A3(new_n639_), .A4(new_n953_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n952_), .A2(new_n959_), .A3(new_n634_), .ZN(new_n960_));
  AND3_X1   g759(.A1(new_n955_), .A2(new_n958_), .A3(new_n960_), .ZN(G1354gat));
  OAI21_X1  g760(.A(KEYINPUT126), .B1(new_n946_), .B2(new_n621_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n904_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  NAND4_X1  g763(.A1(new_n963_), .A2(new_n964_), .A3(new_n655_), .A4(new_n945_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT127), .B(G218gat), .Z(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n962_), .A2(new_n965_), .A3(new_n967_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n956_), .A2(new_n626_), .A3(new_n966_), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1355gat));
endmodule


