//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT10), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G99gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(G106gat), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT9), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n217_), .A2(KEYINPUT64), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n217_), .B2(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n214_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(new_n214_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n211_), .A2(new_n212_), .A3(new_n228_), .ZN(new_n229_));
  NOR4_X1   g028(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n229_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n218_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT67), .ZN(new_n240_));
  OAI22_X1  g039(.A1(new_n235_), .A2(new_n239_), .B1(KEYINPUT8), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n215_), .A2(new_n216_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT8), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n230_), .A2(new_n234_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n242_), .B(new_n244_), .C1(new_n245_), .C2(new_n229_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT68), .B(G71gat), .ZN(new_n248_));
  INV_X1    g047(.A(G78gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n249_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G57gat), .B(G64gat), .Z(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n255_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n227_), .A2(new_n247_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n226_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n219_), .B1(new_n238_), .B2(new_n218_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n220_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n217_), .A2(KEYINPUT64), .A3(new_n220_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n225_), .B1(new_n271_), .B2(new_n214_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n247_), .B1(new_n265_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n260_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT12), .B1(new_n275_), .B2(KEYINPUT69), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n277_), .B(new_n278_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n262_), .B1(new_n275_), .B2(new_n261_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G120gat), .B(G148gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G176gat), .B(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n280_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT71), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n260_), .B1(new_n227_), .B2(new_n247_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n278_), .B1(new_n291_), .B2(new_n277_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n224_), .A2(new_n226_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n293_), .C2(new_n260_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n281_), .B1(new_n295_), .B2(new_n264_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n288_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n288_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n203_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  AOI211_X1 g101(.A(KEYINPUT72), .B(new_n300_), .C1(new_n290_), .C2(new_n298_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n297_), .B1(new_n296_), .B2(new_n288_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n263_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n306_));
  NOR4_X1   g105(.A1(new_n306_), .A2(KEYINPUT71), .A3(new_n281_), .A4(new_n287_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT72), .B1(new_n308_), .B2(new_n300_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n299_), .A2(new_n203_), .A3(new_n301_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT13), .A3(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n304_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G8gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G15gat), .ZN(new_n316_));
  INV_X1    g115(.A(G22gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G15gat), .A2(G22gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G1gat), .A2(G8gat), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n318_), .A2(new_n319_), .B1(KEYINPUT14), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n315_), .B(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(G29gat), .A2(G36gat), .ZN(new_n323_));
  INV_X1    g122(.A(G43gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G29gat), .A2(G36gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G50gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G43gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(G50gat), .B1(new_n332_), .B2(new_n326_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n322_), .B(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G229gat), .A3(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G229gat), .A2(G233gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT78), .Z(new_n338_));
  INV_X1    g137(.A(new_n322_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT15), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n328_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(G50gat), .A3(new_n326_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT15), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(KEYINPUT77), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n341_), .A2(new_n344_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(new_n322_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n322_), .B2(new_n334_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n338_), .B(new_n346_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G113gat), .B(G141gat), .ZN(new_n352_));
  INV_X1    g151(.A(G169gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G197gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n336_), .A2(new_n351_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n336_), .B2(new_n351_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n312_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT99), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT88), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G141gat), .ZN(new_n372_));
  INV_X1    g171(.A(G148gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT89), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT2), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT2), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT3), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n380_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n371_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n372_), .A2(new_n373_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n370_), .B(KEYINPUT1), .Z(new_n385_));
  AOI211_X1 g184(.A(new_n377_), .B(new_n384_), .C1(new_n369_), .C2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389_));
  INV_X1    g188(.A(G113gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n391_), .A2(G120gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G120gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n391_), .B(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(KEYINPUT87), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n388_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n387_), .A2(new_n398_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n366_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT4), .B1(new_n388_), .B2(new_n400_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n365_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n401_), .A2(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n363_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT101), .ZN(new_n410_));
  XOR2_X1   g209(.A(G57gat), .B(G85gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n405_), .A2(new_n407_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT105), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT18), .B(G64gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n428_));
  XOR2_X1   g227(.A(G211gat), .B(G218gat), .Z(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT21), .ZN(new_n431_));
  INV_X1    g230(.A(G204gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G197gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n355_), .A2(G204gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT91), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n434_), .B(KEYINPUT92), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n431_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT93), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n433_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT21), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n430_), .B(new_n436_), .C1(new_n440_), .C2(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n438_), .A2(new_n431_), .A3(new_n430_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT23), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G183gat), .A3(G190gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G183gat), .ZN(new_n453_));
  INV_X1    g252(.A(G190gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT23), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(new_n450_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n452_), .B1(new_n457_), .B2(KEYINPUT84), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G169gat), .A2(G176gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n458_), .A2(KEYINPUT97), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT97), .B1(new_n458_), .B2(new_n463_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT26), .B(G190gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT25), .B(G183gat), .ZN(new_n468_));
  INV_X1    g267(.A(G176gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n353_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n461_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n467_), .A2(new_n468_), .B1(new_n460_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n465_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT22), .B(G169gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n469_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G183gat), .A2(G190gat), .ZN(new_n476_));
  OAI221_X1 g275(.A(new_n475_), .B1(new_n353_), .B2(new_n469_), .C1(new_n456_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n428_), .B1(new_n448_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n439_), .A2(KEYINPUT93), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n442_), .A2(new_n443_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n429_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n446_), .B1(new_n482_), .B2(new_n436_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(KEYINPUT26), .B2(new_n454_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n466_), .B2(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT25), .Z(new_n488_));
  AOI22_X1  g287(.A1(new_n486_), .A2(new_n488_), .B1(KEYINPUT24), .B2(new_n471_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n457_), .C1(KEYINPUT24), .C2(new_n462_), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n458_), .A2(KEYINPUT85), .A3(new_n476_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n458_), .B2(new_n476_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G169gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n353_), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n469_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n470_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n493_), .A2(new_n494_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n483_), .A2(new_n492_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n427_), .B1(new_n479_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n492_), .A2(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n448_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n483_), .A2(new_n477_), .A3(new_n473_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n507_), .A2(KEYINPUT20), .A3(new_n427_), .A4(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n424_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n424_), .A3(new_n509_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT27), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n424_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n479_), .A2(new_n427_), .A3(new_n503_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT103), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(KEYINPUT20), .A3(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n426_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(KEYINPUT103), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n514_), .B1(new_n515_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n513_), .B1(new_n522_), .B2(KEYINPUT27), .ZN(new_n523_));
  XOR2_X1   g322(.A(G78gat), .B(G106gat), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT29), .B1(new_n383_), .B2(new_n386_), .ZN(new_n526_));
  INV_X1    g325(.A(G228gat), .ZN(new_n527_));
  INV_X1    g326(.A(G233gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n448_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n448_), .B2(new_n526_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n387_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G22gat), .B(G50gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT28), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n526_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n529_), .B1(new_n539_), .B2(new_n483_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n448_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n524_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n533_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(KEYINPUT94), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n541_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n525_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT95), .B1(new_n549_), .B2(new_n538_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n546_), .B2(new_n525_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT94), .B(new_n524_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n542_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554_));
  INV_X1    g353(.A(new_n538_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n543_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G15gat), .B(G43gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G227gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT30), .B1(new_n396_), .B2(new_n399_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n394_), .A2(new_n395_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n398_), .A2(KEYINPUT87), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n561_), .A2(new_n492_), .A3(new_n502_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n561_), .A2(new_n565_), .B1(new_n492_), .B2(new_n502_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n560_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G71gat), .B(G99gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n561_), .A2(new_n565_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n506_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n560_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n566_), .A3(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n569_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n572_), .B1(new_n569_), .B2(new_n576_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n557_), .A2(new_n580_), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n543_), .B(new_n579_), .C1(new_n550_), .C2(new_n556_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n420_), .B(new_n523_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n363_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n406_), .A2(new_n365_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n414_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT102), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT102), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n584_), .A2(new_n588_), .A3(new_n414_), .A4(new_n585_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n405_), .A2(KEYINPUT33), .A3(new_n407_), .A4(new_n416_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n514_), .B2(new_n510_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n417_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n511_), .A2(KEYINPUT98), .A3(new_n512_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n591_), .A2(new_n593_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n424_), .A2(KEYINPUT32), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n521_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n505_), .A2(new_n509_), .A3(new_n598_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n521_), .A2(KEYINPUT104), .A3(new_n599_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n602_), .A2(new_n418_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n579_), .A3(new_n557_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n362_), .B1(new_n583_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n293_), .A2(new_n334_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT73), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n293_), .A2(new_n347_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT73), .B1(new_n273_), .B2(new_n345_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(KEYINPUT35), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G134gat), .ZN(new_n618_));
  INV_X1    g417(.A(G162gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT36), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n610_), .B1(new_n293_), .B2(new_n347_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n273_), .A2(KEYINPUT73), .A3(new_n345_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n615_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n628_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n626_), .A2(new_n630_), .A3(new_n631_), .A4(new_n609_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n616_), .A2(new_n623_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT74), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT37), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT75), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n620_), .A2(new_n621_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n623_), .B1(new_n616_), .B2(new_n632_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(new_n633_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT75), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n642_), .A3(KEYINPUT37), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n633_), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n645_), .A2(new_n639_), .B1(new_n621_), .B2(new_n620_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(new_n635_), .B2(KEYINPUT37), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT75), .B(new_n648_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n260_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n339_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT17), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G183gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(G211gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G127gat), .B(G155gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n656_), .B(new_n657_), .Z(new_n658_));
  NOR3_X1   g457(.A1(new_n653_), .A2(new_n654_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(KEYINPUT17), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n653_), .B2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(new_n650_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n608_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(G1gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n420_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT38), .ZN(new_n668_));
  INV_X1    g467(.A(new_n661_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n646_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n608_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G1gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT106), .ZN(G1324gat));
  INV_X1    g474(.A(G8gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n523_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n664_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT107), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n671_), .B2(new_n677_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1325gat));
  AOI21_X1  g484(.A(new_n316_), .B1(new_n671_), .B2(new_n580_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT41), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n664_), .A2(new_n316_), .A3(new_n580_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(new_n557_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n317_), .B1(new_n671_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT42), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n664_), .A2(new_n317_), .A3(new_n690_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n583_), .A2(new_n607_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n646_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n362_), .A2(new_n661_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT108), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n695_), .A2(new_n700_), .A3(new_n697_), .A4(new_n646_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n666_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n644_), .A2(new_n650_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n695_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n705_), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT43), .B(new_n707_), .C1(new_n583_), .C2(new_n607_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n697_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT44), .B(new_n697_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n703_), .B1(new_n714_), .B2(new_n666_), .ZN(G1328gat));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n699_), .A2(new_n716_), .A3(new_n677_), .A4(new_n701_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n711_), .A2(new_n677_), .A3(new_n712_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(KEYINPUT109), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n720_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n722_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n718_), .A2(new_n720_), .A3(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(new_n723_), .ZN(G1329gat));
  NAND4_X1  g526(.A1(new_n711_), .A2(G43gat), .A3(new_n580_), .A4(new_n712_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n699_), .A2(new_n580_), .A3(new_n701_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n324_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(new_n324_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n702_), .B2(new_n690_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n557_), .A2(new_n328_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n713_), .B2(new_n736_), .ZN(G1331gat));
  NOR2_X1   g536(.A1(new_n312_), .A2(new_n361_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n695_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n663_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n666_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n739_), .A2(new_n670_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n666_), .A2(G57gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(G1332gat));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n742_), .B2(new_n677_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT48), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n745_), .A3(new_n677_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n742_), .B2(new_n580_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT49), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n580_), .A2(new_n750_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n740_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1334gat));
  AOI21_X1  g555(.A(new_n249_), .B1(new_n742_), .B2(new_n690_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n740_), .A2(new_n249_), .A3(new_n690_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  NOR3_X1   g559(.A1(new_n312_), .A2(new_n361_), .A3(new_n661_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(KEYINPUT113), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(KEYINPUT113), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT114), .ZN(new_n767_));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n420_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n695_), .A2(new_n646_), .A3(new_n761_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n236_), .A3(new_n666_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1336gat));
  OAI21_X1  g570(.A(G92gat), .B1(new_n767_), .B2(new_n523_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n237_), .A3(new_n677_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1337gat));
  OAI21_X1  g573(.A(G99gat), .B1(new_n766_), .B2(new_n579_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT51), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n579_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n769_), .A2(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n775_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n776_), .A2(KEYINPUT51), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1338gat));
  INV_X1    g581(.A(G106gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n769_), .A2(new_n783_), .A3(new_n690_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n765_), .B(new_n690_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n784_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n784_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795_));
  INV_X1    g594(.A(new_n361_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n304_), .A2(new_n311_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n663_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n304_), .A2(new_n311_), .A3(new_n796_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n799_), .A2(new_n662_), .A3(KEYINPUT54), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n261_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT118), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n295_), .A2(new_n805_), .A3(new_n261_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n262_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n808_));
  NOR2_X1   g607(.A1(new_n306_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT55), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n263_), .B(new_n812_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n287_), .B1(new_n807_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT119), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n361_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n287_), .B(new_n821_), .C1(new_n807_), .C2(new_n814_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n299_), .A2(new_n823_), .A3(new_n361_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n818_), .A2(new_n820_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n335_), .A2(new_n338_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n346_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n826_), .B(new_n356_), .C1(new_n827_), .C2(new_n338_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n358_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT57), .A3(new_n641_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  INV_X1    g634(.A(new_n262_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n805_), .B1(new_n295_), .B2(new_n261_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n261_), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT118), .B(new_n838_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n306_), .A2(new_n811_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n306_), .B2(new_n808_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n288_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n830_), .B1(new_n843_), .B2(new_n816_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n816_), .B(new_n287_), .C1(new_n807_), .C2(new_n814_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n299_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n835_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n829_), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n308_), .B1(new_n843_), .B2(new_n816_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(KEYINPUT58), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n705_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n646_), .B1(new_n825_), .B2(new_n831_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(KEYINPUT57), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n852_), .B2(KEYINPUT57), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n834_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n802_), .B1(new_n856_), .B2(new_n661_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(new_n666_), .A3(new_n582_), .A4(new_n523_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT59), .B1(new_n858_), .B2(KEYINPUT121), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n832_), .A2(new_n641_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n852_), .A2(new_n854_), .A3(KEYINPUT57), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n860_), .A2(new_n863_), .A3(new_n851_), .A4(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n801_), .B1(new_n865_), .B2(new_n669_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(new_n420_), .A3(new_n677_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .A4(new_n582_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n859_), .A2(new_n870_), .A3(G113gat), .A4(new_n361_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n390_), .B1(new_n858_), .B2(new_n796_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1340gat));
  NAND2_X1  g672(.A1(new_n859_), .A2(new_n870_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G120gat), .B1(new_n874_), .B2(new_n312_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n858_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n397_), .B1(new_n312_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n876_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n397_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n874_), .A2(new_n880_), .A3(new_n669_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G127gat), .B1(new_n876_), .B2(new_n661_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n707_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n859_), .A2(new_n870_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n858_), .B2(new_n641_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT122), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n890_), .A3(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n867_), .A2(new_n581_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n796_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n372_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n312_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n373_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n893_), .A2(new_n669_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT123), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n898_), .B(new_n900_), .ZN(G1346gat));
  NOR3_X1   g700(.A1(new_n893_), .A2(new_n619_), .A3(new_n707_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n893_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n646_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n619_), .B2(new_n904_), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n866_), .A2(new_n690_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n677_), .A2(new_n420_), .A3(new_n580_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT62), .B(G169gat), .C1(new_n909_), .C2(new_n796_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n866_), .A2(new_n796_), .A3(new_n690_), .A4(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n474_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n911_), .B2(new_n353_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n910_), .A2(new_n912_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT124), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n910_), .A2(new_n917_), .A3(new_n914_), .A4(new_n912_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1348gat));
  NOR2_X1   g718(.A1(new_n909_), .A2(new_n312_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(G176gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n906_), .B(KEYINPUT125), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n312_), .A3(new_n907_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n923_), .B2(G176gat), .ZN(G1349gat));
  NOR3_X1   g723(.A1(new_n909_), .A2(new_n468_), .A3(new_n669_), .ZN(new_n925_));
  OR3_X1    g724(.A1(new_n922_), .A2(new_n669_), .A3(new_n907_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n453_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n909_), .B2(new_n707_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n646_), .A2(new_n467_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n909_), .B2(new_n929_), .ZN(G1351gat));
  AND2_X1   g729(.A1(new_n581_), .A2(new_n420_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n866_), .A2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n523_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n796_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n355_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n312_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n432_), .ZN(G1353gat));
  INV_X1    g739(.A(new_n936_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n661_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n942_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n942_), .B2(new_n943_), .ZN(G1354gat));
  XNOR2_X1  g745(.A(KEYINPUT127), .B(G218gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n936_), .A2(new_n707_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n941_), .A2(new_n646_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n947_), .ZN(G1355gat));
endmodule


