//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n205_), .A2(new_n210_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n216_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n204_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .A3(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n224_), .A3(new_n212_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n209_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT65), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n208_), .A2(new_n229_), .A3(new_n209_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n215_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n215_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n218_), .A2(new_n219_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n212_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n214_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G36gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G29gat), .ZN(new_n240_));
  INV_X1    g039(.A(G29gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G36gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n240_), .A2(new_n242_), .A3(KEYINPUT69), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT69), .B1(new_n240_), .B2(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n238_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n241_), .A2(G36gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n239_), .A2(G29gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n242_), .A3(KEYINPUT69), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n237_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n245_), .A2(KEYINPUT15), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT15), .B1(new_n245_), .B2(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n236_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n245_), .A2(new_n251_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(new_n214_), .C1(new_n232_), .C2(new_n235_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(new_n258_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n254_), .A2(new_n265_), .A3(new_n259_), .A4(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G134gat), .B(G162gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n267_), .A2(KEYINPUT36), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT37), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n270_), .B(KEYINPUT36), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(KEYINPUT70), .A3(new_n266_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n267_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n271_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n281_), .B2(KEYINPUT37), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n285_));
  XOR2_X1   g084(.A(G71gat), .B(G78gat), .Z(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  INV_X1    g091(.A(G1gat), .ZN(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n290_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n289_), .B(new_n299_), .Z(new_n300_));
  NAND2_X1  g099(.A1(G231gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT17), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(KEYINPUT17), .A3(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n202_), .B1(new_n282_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT5), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n289_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n236_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n289_), .B(new_n214_), .C1(new_n232_), .C2(new_n235_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(KEYINPUT67), .A3(new_n320_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n236_), .A2(KEYINPUT67), .A3(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT64), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n324_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT12), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n236_), .A2(new_n329_), .A3(new_n318_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n236_), .B2(new_n318_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n317_), .B1(new_n326_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n333_), .A3(new_n317_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT13), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n334_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n280_), .A2(new_n277_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n271_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n344_), .A2(new_n272_), .B1(new_n275_), .B2(new_n273_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n311_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT72), .A3(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n312_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G229gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n260_), .A2(new_n299_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n251_), .A2(new_n245_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT73), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n299_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n351_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n349_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(new_n350_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G113gat), .B(G141gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT74), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G169gat), .B(G197gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n354_), .A2(new_n357_), .A3(new_n359_), .A4(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n354_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368_));
  INV_X1    g167(.A(new_n363_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT76), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n364_), .A2(new_n365_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G183gat), .ZN(new_n379_));
  INV_X1    g178(.A(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT23), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G183gat), .A3(G190gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT79), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n382_), .B2(KEYINPUT23), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n381_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G169gat), .ZN(new_n390_));
  INV_X1    g189(.A(G176gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT22), .B(G169gat), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT78), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(KEYINPUT22), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396_));
  AOI21_X1  g195(.A(G176gat), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n392_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  OR3_X1    g197(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n392_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT26), .B(G190gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT77), .B1(new_n379_), .B2(KEYINPUT25), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT25), .B(G183gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n404_), .C1(new_n405_), .C2(KEYINPUT77), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n389_), .A2(new_n398_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(G43gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G15gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT30), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n415_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n412_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT81), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G155gat), .A3(G162gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G141gat), .A2(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n434_), .B2(KEYINPUT82), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AND3_X1   g240(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n434_), .A2(KEYINPUT82), .A3(new_n439_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n427_), .A2(new_n432_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n433_), .A2(new_n438_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT84), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G197gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G204gat), .ZN(new_n453_));
  INV_X1    g252(.A(G204gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G197gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT21), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G211gat), .B(G218gat), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT86), .B1(new_n454_), .B2(G197gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT85), .B1(new_n452_), .B2(G204gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n452_), .A3(G204gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n454_), .A3(G197gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT21), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n459_), .B1(new_n456_), .B2(KEYINPUT21), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n460_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n431_), .B1(new_n427_), .B2(KEYINPUT1), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n437_), .B1(new_n476_), .B2(new_n430_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n440_), .A2(new_n443_), .A3(new_n442_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n447_), .B1(new_n478_), .B2(new_n445_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n475_), .B(KEYINPUT29), .C1(new_n477_), .C2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n451_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n469_), .B1(KEYINPUT21), .B2(new_n467_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT87), .B1(new_n482_), .B2(new_n460_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n470_), .A2(new_n468_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n460_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n433_), .A2(new_n438_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n446_), .A2(new_n448_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT29), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n472_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(KEYINPUT89), .B(new_n422_), .C1(new_n481_), .C2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G22gat), .B(G50gat), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n497_));
  NOR4_X1   g296(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT29), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n496_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n497_), .B1(new_n491_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n449_), .A2(new_n450_), .A3(new_n499_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n495_), .A3(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n488_), .A2(new_n492_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n473_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n451_), .A2(new_n480_), .A3(new_n474_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n422_), .A2(KEYINPUT89), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n494_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n483_), .A2(new_n487_), .B1(new_n491_), .B2(KEYINPUT29), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n508_), .B(new_n422_), .C1(new_n472_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n501_), .A2(new_n504_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n422_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n512_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n422_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n481_), .B2(new_n493_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(new_n514_), .A3(KEYINPUT88), .A4(new_n515_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n511_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n418_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n489_), .A2(new_n490_), .A3(new_n418_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n449_), .A2(KEYINPUT92), .A3(new_n418_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G29gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G85gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT0), .B(G57gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT4), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n491_), .A2(new_n538_), .A3(new_n523_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n530_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n531_), .B(new_n537_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n529_), .A2(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n530_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n544_), .B(new_n535_), .C1(new_n539_), .C2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G8gat), .B(G36gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT18), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G64gat), .B(G92gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n401_), .B1(new_n405_), .B2(new_n403_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n386_), .A2(new_n388_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G169gat), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n392_), .B1(new_n560_), .B2(new_n391_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n383_), .A2(new_n385_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n381_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n563_), .A3(KEYINPUT91), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT91), .B1(new_n561_), .B2(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n559_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n484_), .A2(new_n485_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n556_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n407_), .A2(new_n471_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n555_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT20), .B1(new_n407_), .B2(new_n471_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n551_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n561_), .A2(new_n563_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n578_), .A2(new_n564_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT20), .B1(new_n579_), .B2(new_n471_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n398_), .A2(new_n389_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n402_), .A2(new_n406_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n568_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n554_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n554_), .B1(new_n579_), .B2(new_n471_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n556_), .B1(new_n583_), .B2(new_n568_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n588_), .A3(new_n550_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n543_), .A2(new_n546_), .A3(new_n575_), .A4(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n541_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n529_), .A2(KEYINPUT4), .ZN(new_n592_));
  INV_X1    g391(.A(new_n542_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n535_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT33), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n580_), .A2(new_n584_), .A3(new_n554_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n483_), .A2(new_n487_), .A3(new_n559_), .A4(new_n576_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n555_), .B1(new_n587_), .B2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n585_), .A2(new_n602_), .A3(new_n588_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n551_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n585_), .A2(KEYINPUT93), .A3(new_n588_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n604_), .B2(new_n551_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n539_), .A2(new_n542_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n535_), .B1(new_n609_), .B2(new_n591_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n531_), .B(new_n595_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n606_), .A2(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n522_), .B(KEYINPUT94), .C1(new_n597_), .C2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n518_), .A2(new_n521_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n511_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n571_), .A2(new_n574_), .A3(new_n551_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT27), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n551_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n575_), .A2(new_n589_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n619_), .A2(new_n620_), .B1(new_n621_), .B2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(new_n611_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n613_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n606_), .A2(new_n608_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n623_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n550_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n617_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n611_), .A2(new_n536_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n543_), .A4(new_n546_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT94), .B1(new_n633_), .B2(new_n522_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n421_), .B1(new_n626_), .B2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n622_), .A2(new_n522_), .A3(new_n624_), .A4(new_n420_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n378_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n348_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n293_), .A3(new_n623_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT95), .Z(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT38), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT38), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n281_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n378_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n341_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n311_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n624_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n642_), .A3(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(new_n622_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n348_), .A2(new_n637_), .A3(new_n294_), .A4(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT96), .ZN(new_n652_));
  OAI21_X1  g451(.A(G8gat), .B1(new_n647_), .B2(new_n622_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT98), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT98), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n647_), .B2(new_n421_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n638_), .A2(new_n666_), .A3(new_n420_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  XNOR2_X1  g467(.A(new_n616_), .B(KEYINPUT99), .ZN(new_n669_));
  OAI21_X1  g468(.A(G22gat), .B1(new_n647_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n669_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n638_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1327gat));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n635_), .A2(new_n636_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n282_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT43), .B(new_n345_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n645_), .A2(new_n346_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT101), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n681_), .A2(new_n683_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n623_), .B(new_n684_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G29gat), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n637_), .A2(new_n341_), .A3(new_n311_), .A4(new_n281_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n241_), .A3(new_n623_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT103), .ZN(G1328gat));
  OAI211_X1 g491(.A(new_n650_), .B(new_n684_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n239_), .A3(new_n650_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT45), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1329gat));
  AOI21_X1  g498(.A(G43gat), .B1(new_n689_), .B2(new_n420_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT104), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n420_), .A2(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n704_), .B(new_n705_), .Z(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n689_), .B2(new_n674_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n702_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n616_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  INV_X1    g509(.A(new_n341_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n644_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n712_));
  AND4_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n312_), .A4(new_n347_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n623_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n311_), .B1(new_n377_), .B2(new_n372_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n643_), .A2(new_n711_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n624_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n717_), .B2(new_n622_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n622_), .A2(G64gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT107), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n713_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n717_), .B2(new_n421_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  INV_X1    g527(.A(G71gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n713_), .A2(new_n729_), .A3(new_n420_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n717_), .B2(new_n669_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n713_), .A2(new_n734_), .A3(new_n674_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1335gat));
  AND4_X1   g535(.A1(new_n711_), .A2(new_n712_), .A3(new_n311_), .A4(new_n281_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n623_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT108), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n341_), .A2(new_n644_), .A3(new_n346_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n681_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n624_), .A2(new_n206_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n741_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n737_), .B2(new_n650_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n622_), .A2(new_n207_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT109), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n741_), .B2(new_n746_), .ZN(G1337gat));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n737_), .A2(new_n420_), .A3(new_n203_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n420_), .B(new_n740_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G99gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G99gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT111), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  AND4_X1   g556(.A1(new_n748_), .A2(new_n755_), .A3(KEYINPUT51), .A4(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT112), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n754_), .B2(KEYINPUT111), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n757_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n758_), .A2(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n737_), .A2(new_n204_), .A3(new_n616_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n681_), .A2(new_n616_), .A3(new_n740_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  AND4_X1   g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .A4(G106gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n204_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n767_), .A2(new_n770_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n341_), .A2(new_n716_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n341_), .B2(new_n716_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n345_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n345_), .B(new_n778_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n339_), .A2(new_n334_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n355_), .A2(new_n356_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n349_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n786_), .B2(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n369_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n364_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n784_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n372_), .A2(new_n377_), .A3(new_n336_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n372_), .A2(new_n377_), .A3(KEYINPUT116), .A4(new_n336_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n319_), .A2(KEYINPUT12), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n327_), .B1(new_n799_), .B2(new_n330_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(KEYINPUT55), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n333_), .A2(KEYINPUT117), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(KEYINPUT55), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n320_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n325_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n801_), .A2(new_n803_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n316_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n316_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n792_), .B1(new_n797_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n783_), .B1(new_n813_), .B2(new_n281_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n811_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n316_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n795_), .A2(new_n796_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT57), .B(new_n344_), .C1(new_n819_), .C2(new_n792_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n814_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n790_), .A2(new_n364_), .A3(new_n336_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT58), .B(new_n825_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n282_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n782_), .B1(new_n828_), .B2(new_n311_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NOR4_X1   g630(.A1(new_n650_), .A2(new_n421_), .A3(new_n616_), .A4(new_n624_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n823_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n282_), .B1(new_n834_), .B2(KEYINPUT58), .ZN(new_n835_));
  INV_X1    g634(.A(new_n826_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT119), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n824_), .A2(new_n838_), .A3(new_n282_), .A4(new_n826_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n814_), .A2(new_n837_), .A3(new_n839_), .A4(new_n820_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n311_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n782_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n832_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n833_), .B1(new_n831_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n378_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n847_), .A3(new_n644_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n845_), .B2(new_n341_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n341_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n844_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n845_), .B2(new_n311_), .ZN(new_n855_));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n844_), .A2(new_n856_), .A3(new_n346_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1342gat));
  OAI21_X1  g657(.A(G134gat), .B1(new_n845_), .B2(new_n345_), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n844_), .A2(new_n860_), .A3(new_n281_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1343gat));
  AOI21_X1  g661(.A(new_n782_), .B1(new_n840_), .B2(new_n311_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n421_), .A2(new_n616_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n644_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n711_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n346_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(KEYINPUT120), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(KEYINPUT120), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  NAND2_X1  g674(.A1(new_n865_), .A2(new_n282_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n344_), .A2(G162gat), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n876_), .A2(G162gat), .B1(new_n865_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT121), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n622_), .A2(new_n623_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n420_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n674_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n830_), .A2(new_n880_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n883_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT123), .B1(new_n829_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n560_), .A3(new_n644_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n346_), .B1(new_n821_), .B2(new_n827_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n644_), .B(new_n883_), .C1(new_n889_), .C2(new_n782_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n891_), .B2(new_n390_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n894_), .A3(G169gat), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n888_), .B1(new_n896_), .B2(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n887_), .B2(new_n711_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n863_), .A2(new_n616_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n882_), .A2(new_n391_), .A3(new_n341_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n311_), .A2(new_n405_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n900_), .A2(new_n420_), .A3(new_n346_), .A4(new_n881_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n887_), .A2(new_n903_), .B1(new_n379_), .B2(new_n904_), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n887_), .A2(new_n403_), .A3(new_n281_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n345_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n380_), .B2(new_n907_), .ZN(G1351gat));
  NAND3_X1  g707(.A1(new_n881_), .A2(new_n616_), .A3(new_n421_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n863_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n644_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n452_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(G197gat), .A3(new_n644_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n913_), .A2(KEYINPUT124), .ZN(new_n914_));
  AOI211_X1 g713(.A(new_n912_), .B(new_n914_), .C1(new_n452_), .C2(new_n911_), .ZN(G1352gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n863_), .A2(new_n341_), .A3(new_n909_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n454_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  OAI21_X1  g718(.A(G204gat), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n863_), .A2(KEYINPUT125), .A3(new_n341_), .A4(new_n909_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  INV_X1    g722(.A(new_n909_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n843_), .A2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT125), .B1(new_n925_), .B2(new_n341_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n910_), .A2(new_n919_), .A3(new_n711_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n926_), .A2(new_n916_), .A3(G204gat), .A4(new_n927_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n922_), .A2(new_n923_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n923_), .B1(new_n922_), .B2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1353gat));
  NAND2_X1  g730(.A1(new_n910_), .A2(new_n346_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n932_), .B2(new_n933_), .ZN(G1354gat));
  OR3_X1    g735(.A1(new_n925_), .A2(G218gat), .A3(new_n344_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G218gat), .B1(new_n925_), .B2(new_n345_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1355gat));
endmodule


