//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT83), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT4), .ZN(new_n213_));
  INV_X1    g012(.A(G155gat), .ZN(new_n214_));
  INV_X1    g013(.A(G162gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT84), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT87), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT87), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT3), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n225_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT88), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n221_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G141gat), .ZN(new_n237_));
  INV_X1    g036(.A(G148gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n219_), .B2(KEYINPUT1), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n244_), .A2(KEYINPUT85), .A3(G155gat), .A4(G162gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n216_), .A2(new_n247_), .A3(new_n218_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n236_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n213_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT97), .B(new_n212_), .C1(new_n250_), .C2(KEYINPUT98), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT97), .ZN(new_n257_));
  INV_X1    g056(.A(new_n232_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(new_n230_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n234_), .B(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n261_), .A3(new_n225_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n246_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n248_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n262_), .A2(new_n221_), .B1(new_n265_), .B2(new_n241_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT98), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n236_), .A2(new_n257_), .A3(new_n249_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n211_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n208_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n256_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT99), .A3(KEYINPUT4), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT99), .B1(new_n274_), .B2(KEYINPUT4), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n255_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n252_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G57gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n279_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT102), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n274_), .A2(KEYINPUT4), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT99), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n254_), .B1(new_n289_), .B2(new_n275_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n279_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT102), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n278_), .A2(new_n293_), .A3(new_n279_), .A4(new_n283_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n285_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n296_), .A2(KEYINPUT24), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT23), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n305_), .B2(new_n303_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n305_), .B2(new_n303_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G169gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT30), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G71gat), .B(G99gat), .ZN(new_n319_));
  INV_X1    g118(.A(G43gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(G15gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n316_), .A2(new_n317_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n272_), .B(KEYINPUT31), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT22), .B(G169gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT96), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n311_), .A2(new_n297_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n301_), .A2(KEYINPUT95), .A3(new_n307_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT95), .B1(new_n301_), .B2(new_n307_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G197gat), .ZN(new_n355_));
  INV_X1    g154(.A(G197gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G204gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G218gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G211gat), .ZN(new_n360_));
  INV_X1    g159(.A(G211gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G218gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(KEYINPUT21), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n358_), .A2(new_n363_), .A3(new_n366_), .A4(KEYINPUT21), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT21), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n355_), .A2(new_n357_), .A3(KEYINPUT91), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n356_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT21), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n368_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n343_), .B1(new_n353_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n355_), .A2(new_n357_), .A3(KEYINPUT91), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT21), .B1(new_n355_), .B2(KEYINPUT91), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n360_), .B(new_n362_), .C1(new_n358_), .C2(KEYINPUT21), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT92), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n371_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n384_), .A2(new_n385_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n314_), .A3(new_n308_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n342_), .B1(new_n379_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n308_), .A2(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n390_), .A2(new_n350_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n386_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n343_), .B1(new_n378_), .B2(new_n315_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n392_), .A2(new_n342_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n339_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n387_), .B(KEYINPUT20), .C1(new_n391_), .C2(new_n386_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n341_), .B1(new_n391_), .B2(new_n386_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n396_), .A2(new_n341_), .B1(new_n397_), .B2(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n338_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n396_), .A2(new_n341_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n386_), .A2(new_n349_), .A3(new_n308_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n342_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n339_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n398_), .B2(new_n338_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n400_), .A2(new_n401_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n334_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n266_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT28), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n236_), .B2(new_n249_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT90), .B1(new_n386_), .B2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n224_), .B1(new_n418_), .B2(new_n258_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n220_), .B1(new_n419_), .B2(new_n261_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n249_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT29), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n378_), .ZN(new_n424_));
  INV_X1    g223(.A(G78gat), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n417_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n417_), .B2(new_n424_), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n386_), .A2(new_n416_), .A3(KEYINPUT90), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n423_), .B1(new_n422_), .B2(new_n378_), .ZN(new_n431_));
  OAI21_X1  g230(.A(G78gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n417_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n433_));
  AOI21_X1  g232(.A(G106gat), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n415_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n428_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(G106gat), .A3(new_n433_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(G228gat), .A4(G233gat), .ZN(new_n439_));
  AND4_X1   g238(.A1(KEYINPUT89), .A2(new_n435_), .A3(new_n436_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n438_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(new_n415_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n443_), .B2(new_n439_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n414_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n435_), .A2(KEYINPUT89), .A3(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT94), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n413_), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n295_), .B(new_n408_), .C1(new_n445_), .C2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n407_), .A2(new_n285_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n334_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n445_), .A2(new_n449_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n289_), .A2(new_n275_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n283_), .B1(new_n274_), .B2(new_n253_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n400_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n291_), .B1(new_n456_), .B2(new_n255_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n283_), .ZN(new_n464_));
  NOR4_X1   g263(.A1(new_n290_), .A2(KEYINPUT33), .A3(new_n291_), .A4(new_n286_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n461_), .B(KEYINPUT101), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n402_), .A2(new_n404_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n398_), .B2(new_n468_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n295_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n455_), .A2(new_n466_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n450_), .B1(new_n454_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT65), .Z(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G85gat), .A3(G92gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT10), .B(G99gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G85gat), .B(G92gat), .ZN(new_n486_));
  OAI221_X1 g285(.A(new_n484_), .B1(new_n485_), .B2(G106gat), .C1(new_n483_), .C2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT8), .ZN(new_n489_));
  INV_X1    g288(.A(new_n486_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n489_), .B(new_n490_), .C1(new_n482_), .C2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n481_), .A2(KEYINPUT67), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n481_), .A2(KEYINPUT67), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n497_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT8), .B1(new_n499_), .B2(new_n486_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n488_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G29gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT70), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n502_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT15), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n505_), .A2(new_n509_), .A3(KEYINPUT15), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n501_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n501_), .A2(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT34), .Z(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n516_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n520_), .B(KEYINPUT73), .Z(new_n523_));
  AND2_X1   g322(.A1(new_n518_), .A2(new_n519_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT74), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n527_), .B(new_n528_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n521_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G190gat), .B(G218gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT72), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n521_), .B(new_n538_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT16), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n549_));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT68), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555_));
  INV_X1    g354(.A(G1gat), .ZN(new_n556_));
  INV_X1    g355(.A(G8gat), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G8gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n546_), .B1(new_n554_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n554_), .B2(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n553_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n567_), .A2(new_n545_), .A3(new_n544_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n566_), .B2(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n476_), .A2(new_n540_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n501_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n554_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT64), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n501_), .A2(new_n554_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n577_), .A2(KEYINPUT12), .A3(new_n566_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n584_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n583_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n576_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n586_), .A2(new_n589_), .A3(new_n576_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT79), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n510_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n561_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n505_), .A2(new_n509_), .A3(KEYINPUT79), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n606_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT80), .B1(new_n608_), .B2(new_n561_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT80), .ZN(new_n610_));
  AOI211_X1 g409(.A(new_n610_), .B(new_n605_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n602_), .B(new_n607_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n606_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT79), .B1(new_n505_), .B2(new_n509_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n561_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n610_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n608_), .A2(KEYINPUT80), .A3(new_n561_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n605_), .B2(new_n514_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n612_), .B(new_n616_), .C1(new_n622_), .C2(new_n602_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n612_), .B1(new_n622_), .B2(new_n602_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n615_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n624_), .B2(new_n615_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n601_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n571_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n295_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT103), .Z(new_n634_));
  INV_X1    g433(.A(new_n623_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n624_), .A2(new_n615_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT81), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n624_), .A2(new_n625_), .A3(new_n615_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n476_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n516_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n501_), .A2(new_n514_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n525_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n527_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n522_), .A2(KEYINPUT74), .A3(new_n525_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n522_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n644_), .A2(new_n645_), .B1(new_n646_), .B2(new_n520_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n534_), .B(KEYINPUT75), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n539_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT37), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT76), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT76), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n652_), .A3(KEYINPUT37), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n655_));
  INV_X1    g454(.A(new_n534_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n539_), .B(new_n655_), .C1(new_n647_), .C2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT78), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT78), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n535_), .A2(new_n659_), .A3(new_n539_), .A4(new_n655_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n570_), .B1(new_n654_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n601_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n640_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n556_), .A3(new_n295_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT38), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n634_), .A2(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(new_n407_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n557_), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n571_), .A2(new_n630_), .A3(new_n671_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G8gat), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT39), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT39), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g477(.A1(new_n666_), .A2(G15gat), .A3(new_n453_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT104), .Z(new_n680_));
  OAI21_X1  g479(.A(G15gat), .B1(new_n631_), .B2(new_n453_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n682_), .A3(new_n683_), .ZN(G1326gat));
  OAI21_X1  g483(.A(G22gat), .B1(new_n631_), .B2(new_n455_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n455_), .A2(G22gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT105), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n666_), .B2(new_n688_), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n540_), .A2(new_n570_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n664_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n640_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n295_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n570_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n652_), .B1(new_n649_), .B2(KEYINPUT37), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n649_), .A2(new_n652_), .A3(KEYINPUT37), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n661_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n408_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n455_), .A2(new_n632_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n474_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n447_), .A2(new_n448_), .A3(new_n413_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n413_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n452_), .A2(new_n453_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n701_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  INV_X1    g508(.A(new_n698_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n629_), .B(new_n695_), .C1(new_n699_), .C2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT106), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n453_), .B(new_n452_), .C1(new_n702_), .C2(new_n705_), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT43), .B(new_n698_), .C1(new_n715_), .C2(new_n701_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n630_), .B(new_n570_), .C1(new_n714_), .C2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n713_), .A2(new_n720_), .B1(KEYINPUT44), .B2(new_n712_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n295_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n694_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n692_), .A2(G36gat), .A3(new_n407_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n671_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n713_), .B2(new_n720_), .ZN(new_n728_));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n726_), .B(KEYINPUT46), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  NAND2_X1  g533(.A1(new_n712_), .A2(KEYINPUT44), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n453_), .A2(new_n320_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n718_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n735_), .B(new_n736_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n320_), .B1(new_n692_), .B2(new_n453_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  OR3_X1    g544(.A1(new_n692_), .A2(G50gat), .A3(new_n455_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n705_), .B(new_n735_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G50gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G50gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1331gat));
  NOR2_X1   g550(.A1(new_n601_), .A2(new_n628_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n571_), .A2(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT109), .Z(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G57gat), .B1(new_n755_), .B2(new_n632_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n708_), .A2(new_n752_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n663_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n632_), .A2(G57gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n762_), .A3(new_n671_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n754_), .A2(new_n671_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G64gat), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT48), .B(new_n762_), .C1(new_n754_), .C2(new_n671_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n769_), .A3(new_n334_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n754_), .A2(new_n334_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G71gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT49), .B(new_n769_), .C1(new_n754_), .C2(new_n334_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1334gat));
  NAND3_X1  g574(.A1(new_n758_), .A2(new_n425_), .A3(new_n705_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n754_), .A2(new_n705_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(G78gat), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT50), .B(new_n425_), .C1(new_n754_), .C2(new_n705_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n699_), .A2(new_n711_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n570_), .A3(new_n752_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n632_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n757_), .A2(new_n690_), .ZN(new_n785_));
  INV_X1    g584(.A(G85gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n295_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1336gat));
  AOI21_X1  g587(.A(G92gat), .B1(new_n785_), .B2(new_n671_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n783_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n671_), .A2(G92gat), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT110), .Z(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n790_), .B2(new_n792_), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n783_), .B2(new_n453_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n453_), .A2(new_n485_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT111), .B1(new_n785_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n797_), .B(new_n798_), .Z(G1338gat));
  NAND3_X1  g598(.A1(new_n785_), .A2(new_n428_), .A3(new_n705_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n782_), .A2(new_n705_), .A3(new_n570_), .A4(new_n752_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n698_), .A2(new_n639_), .A3(new_n601_), .A4(new_n695_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n662_), .A2(new_n639_), .A3(new_n601_), .A4(new_n809_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n622_), .A2(new_n602_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n607_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n616_), .C1(new_n817_), .C2(new_n602_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n597_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n628_), .A2(new_n593_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n586_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n585_), .A2(new_n584_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(KEYINPUT55), .A3(new_n583_), .A4(new_n581_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n585_), .A2(new_n584_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT12), .B1(new_n577_), .B2(new_n578_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n588_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n825_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n575_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n821_), .A2(KEYINPUT114), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n628_), .A2(new_n835_), .A3(new_n593_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n820_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n814_), .B1(new_n837_), .B2(new_n540_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n833_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n593_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT114), .B1(new_n639_), .B2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n841_), .A3(new_n836_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n820_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n540_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT57), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n575_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n593_), .B(new_n818_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n846_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n850_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n839_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n851_), .A2(new_n854_), .A3(new_n654_), .A4(new_n661_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n838_), .A2(new_n845_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n813_), .B1(new_n856_), .B2(new_n570_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n455_), .A2(new_n295_), .A3(new_n700_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n807_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n837_), .A2(new_n814_), .A3(new_n540_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n570_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n811_), .A2(new_n812_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n858_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(KEYINPUT116), .A3(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n859_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n628_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n858_), .B(new_n871_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT118), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n873_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n864_), .A2(new_n865_), .A3(new_n870_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n639_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n869_), .B1(new_n882_), .B2(new_n868_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n867_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n874_), .A2(new_n875_), .A3(new_n601_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n884_), .B2(new_n887_), .ZN(G1341gat));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889_));
  INV_X1    g688(.A(G127gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n570_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n859_), .A2(new_n866_), .A3(new_n695_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n894_), .A2(new_n890_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n889_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n880_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n891_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n890_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(KEYINPUT119), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n901_), .ZN(G1342gat));
  AOI21_X1  g701(.A(G134gat), .B1(new_n867_), .B2(new_n540_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n876_), .A2(new_n881_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n710_), .A2(G134gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT120), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n455_), .A2(new_n334_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n295_), .A3(new_n407_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT121), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n864_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n628_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n664_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n695_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  INV_X1    g717(.A(new_n911_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G162gat), .B1(new_n919_), .B2(new_n698_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n911_), .A2(new_n215_), .A3(new_n540_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n295_), .A2(new_n407_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n705_), .A2(new_n453_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n628_), .A4(new_n927_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n928_), .A2(G169gat), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n927_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n931_), .B2(new_n639_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n929_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n930_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n628_), .A2(new_n345_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT123), .Z(new_n936_));
  OAI22_X1  g735(.A1(new_n933_), .A2(new_n934_), .B1(new_n931_), .B2(new_n936_), .ZN(G1348gat));
  NOR2_X1   g736(.A1(new_n931_), .A2(new_n601_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n346_), .ZN(G1349gat));
  NOR2_X1   g738(.A1(new_n931_), .A2(new_n570_), .ZN(new_n940_));
  MUX2_X1   g739(.A(G183gat), .B(new_n299_), .S(new_n940_), .Z(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n931_), .B2(new_n698_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n540_), .A2(new_n300_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n931_), .B2(new_n943_), .ZN(G1351gat));
  XOR2_X1   g743(.A(KEYINPUT124), .B(G197gat), .Z(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n925_), .A2(new_n908_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n639_), .ZN(new_n948_));
  MUX2_X1   g747(.A(new_n945_), .B(new_n946_), .S(new_n948_), .Z(G1352gat));
  INV_X1    g748(.A(new_n947_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n664_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(G204gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(G204gat), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n951_), .B2(new_n954_), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n925_), .A2(new_n695_), .A3(new_n908_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT63), .B(G211gat), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  AND3_X1   g759(.A1(new_n956_), .A2(new_n959_), .A3(new_n960_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n956_), .B2(new_n960_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n958_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n958_), .B(KEYINPUT127), .C1(new_n961_), .C2(new_n962_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n947_), .B2(new_n698_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n540_), .A2(new_n359_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n947_), .B2(new_n969_), .ZN(G1355gat));
endmodule


