//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n206_));
  INV_X1    g005(.A(G155gat), .ZN(new_n207_));
  INV_X1    g006(.A(G162gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT1), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n211_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G155gat), .A3(G162gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT87), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n202_), .B(new_n205_), .C1(new_n217_), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n202_), .B1(new_n222_), .B2(KEYINPUT88), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT88), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n202_), .A2(KEYINPUT88), .A3(new_n222_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n209_), .A2(new_n210_), .B1(G155gat), .B2(G162gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT89), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n233_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(KEYINPUT2), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n226_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n227_), .ZN(new_n237_));
  OAI211_X1 g036(.A(KEYINPUT89), .B(new_n231_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n221_), .B1(new_n232_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G113gat), .B(G120gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n248_), .A3(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n246_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n249_), .B(new_n250_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G57gat), .B(G85gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n216_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n261_), .A2(new_n214_), .B1(new_n210_), .B2(new_n209_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n219_), .B(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n262_), .A2(new_n264_), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n231_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n265_), .A2(new_n205_), .B1(new_n268_), .B2(new_n238_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G22gat), .B(G50gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n240_), .A2(KEYINPUT29), .A3(new_n272_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n240_), .A2(KEYINPUT29), .ZN(new_n284_));
  OR2_X1    g083(.A1(G211gat), .A2(G218gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G211gat), .A2(G218gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT92), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n285_), .A2(new_n289_), .A3(new_n286_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n288_), .A2(new_n290_), .B1(new_n292_), .B2(KEYINPUT21), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT21), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n291_), .B(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n283_), .B1(new_n284_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n291_), .A2(new_n297_), .ZN(new_n301_));
  INV_X1    g100(.A(G197gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(G204gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(G204gat), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT21), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n288_), .B(new_n290_), .C1(new_n301_), .C2(new_n305_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n294_), .A2(new_n295_), .B1(new_n297_), .B2(new_n291_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n283_), .ZN(new_n309_));
  AOI211_X1 g108(.A(new_n308_), .B(new_n309_), .C1(new_n240_), .C2(KEYINPUT29), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n282_), .B1(new_n300_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n284_), .A2(new_n299_), .A3(new_n283_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n268_), .A2(new_n238_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n270_), .B1(new_n313_), .B2(new_n221_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n314_), .B2(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n315_), .A3(new_n281_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(KEYINPUT91), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT93), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT93), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n311_), .A2(new_n319_), .A3(new_n316_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n280_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n317_), .A2(KEYINPUT93), .B1(new_n279_), .B2(new_n278_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n260_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT82), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(new_n325_), .A3(G183gat), .A4(G190gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G183gat), .ZN(new_n333_));
  INV_X1    g132(.A(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n324_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT96), .B1(new_n343_), .B2(new_n338_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(new_n324_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n329_), .A2(new_n326_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n352_), .B2(KEYINPUT95), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n329_), .A2(new_n326_), .B1(new_n350_), .B2(new_n349_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  AND2_X1   g154(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n354_), .A2(new_n355_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n336_), .A2(new_n345_), .B1(new_n353_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT97), .B1(new_n361_), .B2(new_n308_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n353_), .A2(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n332_), .A2(new_n335_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n345_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n299_), .ZN(new_n369_));
  AND2_X1   g168(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n357_), .A2(new_n356_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n373_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n365_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n346_), .B2(new_n324_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .A4(KEYINPUT81), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n332_), .A4(new_n351_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n329_), .A2(new_n326_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n383_), .A2(new_n365_), .A3(new_n384_), .A4(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n386_), .A3(new_n308_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n362_), .A2(new_n369_), .A3(KEYINPUT20), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT19), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT94), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n361_), .B2(new_n308_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n390_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n380_), .A2(new_n332_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n377_), .A2(new_n378_), .B1(new_n350_), .B2(new_n349_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n365_), .B1(new_n382_), .B2(KEYINPUT83), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n348_), .A2(KEYINPUT83), .A3(new_n335_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n397_), .A2(new_n398_), .B1(new_n401_), .B2(new_n384_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n395_), .B(new_n396_), .C1(new_n402_), .C2(new_n308_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT18), .B(G64gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n393_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT27), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n388_), .A2(new_n392_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT102), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n367_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n361_), .A2(KEYINPUT102), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n308_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n417_));
  NAND2_X1  g216(.A1(new_n381_), .A2(new_n386_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n299_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n396_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n407_), .B1(new_n412_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT103), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n393_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT103), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n424_), .B(new_n407_), .C1(new_n412_), .C2(new_n420_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n411_), .B1(new_n426_), .B2(KEYINPUT27), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT104), .B1(new_n323_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n322_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n311_), .A2(new_n319_), .A3(new_n316_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(KEYINPUT93), .B2(new_n317_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n431_), .B2(new_n280_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n423_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n363_), .A2(new_n366_), .A3(KEYINPUT102), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT102), .B1(new_n363_), .B2(new_n366_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n299_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n417_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n402_), .B2(new_n308_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n390_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n394_), .B1(new_n402_), .B2(new_n308_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(new_n391_), .A3(new_n362_), .A4(new_n369_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n424_), .B1(new_n442_), .B2(new_n407_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT27), .B1(new_n433_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n411_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT104), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n432_), .A2(new_n446_), .A3(new_n447_), .A4(new_n260_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT100), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n393_), .A3(new_n403_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n442_), .A2(new_n449_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n451_), .B(new_n452_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n257_), .B1(KEYINPUT99), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(KEYINPUT99), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n247_), .A2(new_n251_), .A3(new_n256_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n409_), .A2(new_n410_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n245_), .A2(new_n250_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n256_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n249_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n460_), .B(new_n461_), .C1(new_n462_), .C2(new_n250_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n454_), .A2(KEYINPUT99), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n459_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n453_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n321_), .A2(new_n322_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n428_), .A2(new_n448_), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n402_), .B(KEYINPUT30), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(G71gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n243_), .B(KEYINPUT31), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT84), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G227gat), .A2(G233gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  OR2_X1    g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n476_), .A2(new_n480_), .A3(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n469_), .A2(KEYINPUT105), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT105), .B1(new_n469_), .B2(new_n484_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n260_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n467_), .A2(new_n446_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n485_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT72), .B(G22gat), .ZN(new_n492_));
  INV_X1    g291(.A(G15gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G1gat), .ZN(new_n495_));
  INV_X1    g294(.A(G8gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G8gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n500_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT77), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G229gat), .A3(G233gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT78), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n503_), .B(KEYINPUT15), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n500_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n500_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n503_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT79), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT78), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n505_), .A2(new_n515_), .A3(G229gat), .A4(G233gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n507_), .A2(new_n514_), .A3(new_n516_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G71gat), .B(G78gat), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n529_), .A3(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT6), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n535_));
  OR3_X1    g334(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  XOR2_X1   g337(.A(G85gat), .B(G92gat), .Z(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT67), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT10), .B(G99gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(G106gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT65), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G85gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT9), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(G85gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(G92gat), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n539_), .A2(KEYINPUT9), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n549_), .A2(new_n554_), .A3(new_n534_), .A4(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n532_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT64), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n556_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n544_), .B2(new_n540_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n532_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n532_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT12), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n558_), .A2(new_n561_), .A3(new_n564_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(KEYINPUT66), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT66), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n571_), .A3(new_n532_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n565_), .A2(new_n566_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n569_), .B1(new_n575_), .B2(new_n561_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G204gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT5), .B(G176gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n576_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(KEYINPUT68), .B2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n491_), .A2(new_n525_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n547_), .A2(new_n556_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n590_), .A2(new_n508_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n563_), .A2(new_n503_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT69), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n591_), .B(new_n594_), .C1(new_n596_), .C2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n208_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT70), .B(G134gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT36), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT73), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n500_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n566_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT17), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT17), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n621_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT75), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n621_), .A2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n632_), .B2(KEYINPUT75), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT76), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n617_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n589_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n637_), .A2(G1gat), .A3(new_n260_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n589_), .A2(new_n609_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n260_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1324gat));
  OAI21_X1  g443(.A(G8gat), .B1(new_n642_), .B2(new_n446_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n589_), .A2(new_n496_), .A3(new_n427_), .A4(new_n636_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n642_), .B2(new_n484_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT41), .Z(new_n651_));
  NOR3_X1   g450(.A1(new_n637_), .A2(G15gat), .A3(new_n484_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT107), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1326gat));
  XNOR2_X1  g453(.A(new_n467_), .B(KEYINPUT108), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G22gat), .B1(new_n642_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n637_), .B2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n469_), .A2(new_n484_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n488_), .A2(new_n489_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n469_), .A2(KEYINPUT105), .A3(new_n484_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n617_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT43), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT109), .B(new_n671_), .C1(new_n667_), .C2(new_n617_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n635_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n588_), .A3(new_n525_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n661_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n617_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n669_), .B1(new_n491_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n671_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n668_), .A2(new_n669_), .A3(KEYINPUT43), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n677_), .A2(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n684_), .A2(KEYINPUT110), .A3(new_n260_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT110), .B1(new_n684_), .B2(new_n260_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(G29gat), .A3(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n491_), .A2(new_n609_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n675_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n260_), .A2(G29gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  OAI21_X1  g490(.A(G36gat), .B1(new_n684_), .B2(new_n446_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n689_), .A2(G36gat), .A3(new_n446_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT45), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1329gat));
  INV_X1    g496(.A(new_n689_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G43gat), .B1(new_n698_), .B2(new_n487_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n677_), .A2(new_n683_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n487_), .A2(G43gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n704_), .A3(new_n655_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n700_), .A2(new_n432_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G50gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT111), .B(new_n704_), .C1(new_n700_), .C2(new_n432_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n491_), .A2(new_n635_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n587_), .A2(new_n524_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n609_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n260_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT113), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n678_), .A3(new_n712_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n260_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n716_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n713_), .B2(new_n446_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n446_), .A2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n717_), .B2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT114), .Z(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n713_), .B2(new_n484_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n484_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n717_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n713_), .B2(new_n656_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n656_), .A2(G78gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n717_), .B2(new_n734_), .ZN(G1335gat));
  NAND2_X1  g534(.A1(new_n712_), .A2(new_n635_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n688_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n260_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n673_), .A2(new_n736_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n553_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n260_), .B1(new_n743_), .B2(new_n551_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n742_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n739_), .B2(new_n427_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n427_), .A2(G92gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  NOR3_X1   g547(.A1(new_n738_), .A2(new_n548_), .A3(new_n484_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(new_n487_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G99gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  OAI211_X1 g552(.A(new_n432_), .B(new_n737_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n682_), .A2(KEYINPUT116), .A3(new_n432_), .A4(new_n737_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n756_), .A2(new_n757_), .A3(new_n760_), .A4(G106gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n738_), .A2(G106gat), .A3(new_n467_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n569_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n558_), .A2(new_n573_), .A3(new_n568_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n560_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n567_), .B1(new_n557_), .B2(KEYINPUT12), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n561_), .A4(new_n564_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n580_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT118), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n779_), .A3(new_n580_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT119), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n777_), .A2(new_n784_), .A3(new_n778_), .A4(new_n780_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n576_), .A2(new_n580_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n505_), .A2(new_n513_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n513_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n511_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n520_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n794_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n523_), .A3(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n581_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n609_), .C1(new_n789_), .C2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n786_), .A2(new_n788_), .B1(new_n581_), .B2(new_n797_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n610_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n787_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n776_), .A2(new_n778_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n783_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n797_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n807_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n617_), .A3(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n799_), .A2(new_n802_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n634_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n636_), .A2(new_n525_), .A3(new_n587_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n484_), .A2(new_n489_), .A3(new_n260_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n524_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(new_n635_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n815_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n817_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n524_), .A2(G113gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n820_), .B1(new_n827_), .B2(new_n828_), .ZN(G1340gat));
  XNOR2_X1  g628(.A(KEYINPUT121), .B(G120gat), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT122), .Z(new_n833_));
  OAI211_X1 g632(.A(new_n819_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT124), .B1(new_n826_), .B2(new_n587_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n821_), .A2(new_n838_), .A3(new_n588_), .A4(new_n825_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n830_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n819_), .B2(new_n674_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n641_), .A2(G127gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n827_), .B2(new_n843_), .ZN(G1342gat));
  AOI21_X1  g643(.A(G134gat), .B1(new_n819_), .B2(new_n610_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n617_), .A2(G134gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n827_), .B2(new_n846_), .ZN(G1343gat));
  AOI21_X1  g646(.A(new_n487_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n848_), .A2(new_n740_), .A3(new_n446_), .A4(new_n432_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n525_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n587_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n204_), .ZN(G1345gat));
  NOR2_X1   g652(.A1(new_n849_), .A2(new_n635_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT61), .B(G155gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  NOR3_X1   g655(.A1(new_n849_), .A2(new_n208_), .A3(new_n678_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n208_), .B1(new_n849_), .B2(new_n609_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT125), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(KEYINPUT125), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n488_), .A2(new_n446_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n823_), .A2(new_n524_), .A3(new_n656_), .A4(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G169gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n655_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n342_), .A2(new_n344_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n866_), .A2(new_n524_), .A3(new_n867_), .A4(new_n863_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT62), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT62), .B1(new_n864_), .B2(G169gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n862_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(KEYINPUT126), .A3(new_n871_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1348gat));
  NAND2_X1  g676(.A1(new_n816_), .A2(new_n467_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(G176gat), .A3(new_n588_), .A4(new_n863_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n866_), .A2(new_n863_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n337_), .B1(new_n881_), .B2(new_n587_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n881_), .A2(new_n358_), .A3(new_n634_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n879_), .A2(new_n674_), .A3(new_n863_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n333_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n881_), .B2(new_n678_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n610_), .A2(new_n359_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n881_), .B2(new_n888_), .ZN(G1351gat));
  AND2_X1   g688(.A1(new_n848_), .A2(new_n427_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n323_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n525_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n302_), .ZN(G1352gat));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT127), .B(G204gat), .Z(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n588_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n892_), .A2(new_n587_), .B1(new_n898_), .B2(G204gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1353gat));
  XNOR2_X1  g699(.A(KEYINPUT63), .B(G211gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n895_), .A2(new_n641_), .A3(new_n901_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n892_), .A2(new_n634_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1354gat));
  AND3_X1   g703(.A1(new_n895_), .A2(G218gat), .A3(new_n617_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G218gat), .B1(new_n895_), .B2(new_n610_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


