//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT84), .B1(new_n204_), .B2(new_n205_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n202_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n204_), .A2(new_n205_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n210_), .A2(new_n212_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(G228gat), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G78gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n225_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT21), .ZN(new_n239_));
  INV_X1    g038(.A(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n234_), .B1(new_n240_), .B2(KEYINPUT87), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n240_), .B2(new_n234_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n239_), .B1(KEYINPUT21), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n222_), .B2(new_n221_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G22gat), .B(G50gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n233_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n233_), .A2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT76), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT76), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(G183gat), .A3(G190gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT23), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT79), .ZN(new_n259_));
  AND2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .A4(KEYINPUT23), .ZN(new_n264_));
  OR2_X1    g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n267_), .B2(KEYINPUT22), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT78), .A3(G169gat), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n271_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n267_), .A2(KEYINPUT77), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n267_), .A2(KEYINPUT77), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT22), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n269_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n280_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n269_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n260_), .A2(new_n261_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT23), .B1(new_n255_), .B2(new_n257_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n284_), .B(new_n285_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n279_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT80), .ZN(new_n290_));
  INV_X1    g089(.A(new_n243_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n279_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n265_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n269_), .B1(new_n297_), .B2(new_n268_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n284_), .A2(new_n263_), .A3(new_n285_), .A4(new_n264_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n295_), .B1(new_n243_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n253_), .B1(new_n294_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n243_), .B2(new_n301_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n279_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n292_), .B1(new_n279_), .B2(new_n288_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n243_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT88), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT88), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n243_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n304_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n303_), .B1(new_n311_), .B2(new_n253_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G8gat), .B(G36gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  AOI211_X1 g118(.A(new_n252_), .B(new_n304_), .C1(new_n308_), .C2(new_n310_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n303_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n304_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n290_), .A2(new_n293_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n309_), .B1(new_n327_), .B2(new_n243_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n310_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT92), .A3(new_n252_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n302_), .B(new_n253_), .C1(new_n327_), .C2(new_n243_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT92), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n311_), .B2(new_n253_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n317_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n325_), .B1(new_n335_), .B2(KEYINPUT96), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT96), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n337_), .B(new_n317_), .C1(new_n331_), .C2(new_n334_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n324_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT97), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT97), .B(new_n324_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n250_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G43gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G15gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n345_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n327_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n327_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT82), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n353_), .A2(new_n349_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G127gat), .B(G134gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n361_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT83), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT31), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n359_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT91), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  INV_X1    g180(.A(new_n364_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n363_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI22_X1  g183(.A1(new_n384_), .A2(new_n366_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n209_), .A2(new_n214_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n202_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n216_), .A2(new_n219_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n362_), .A2(new_n364_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n381_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n389_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT4), .B1(new_n393_), .B2(new_n368_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n392_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n380_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n385_), .A2(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT4), .ZN(new_n401_));
  INV_X1    g200(.A(new_n394_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n397_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n377_), .B(new_n378_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n398_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n406_), .A3(KEYINPUT93), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n380_), .C1(new_n396_), .C2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT95), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n373_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n370_), .A2(new_n372_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n312_), .B2(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n330_), .A2(new_n252_), .B1(KEYINPUT92), .B2(new_n332_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n311_), .A2(new_n418_), .A3(new_n253_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT32), .B(new_n317_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n414_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n399_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n404_), .B1(new_n400_), .B2(new_n395_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT33), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n423_), .B1(new_n399_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n249_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n421_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n416_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n413_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n250_), .B1(new_n339_), .B2(new_n411_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n343_), .A2(new_n412_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G57gat), .B(G64gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT11), .ZN(new_n436_));
  XOR2_X1   g235(.A(G71gat), .B(G78gat), .Z(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n435_), .A2(KEYINPUT11), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G85gat), .B(G92gat), .Z(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT10), .B(G99gat), .Z(new_n442_));
  AOI22_X1  g241(.A1(KEYINPUT9), .A2(new_n441_), .B1(new_n442_), .B2(new_n231_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT6), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n443_), .B(new_n445_), .C1(KEYINPUT9), .C2(new_n446_), .ZN(new_n447_));
  OR4_X1    g246(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n231_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT7), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n441_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT8), .B1(new_n441_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n447_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n454_), .A2(new_n456_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n438_), .B(new_n440_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n460_), .A2(KEYINPUT12), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n458_), .A2(new_n459_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n440_), .A2(new_n438_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT12), .A3(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n464_), .B2(new_n460_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G120gat), .B(G148gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT5), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G176gat), .B(G204gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n471_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n469_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n477_), .B1(new_n480_), .B2(new_n472_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(KEYINPUT68), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n483_), .B(new_n477_), .C1(new_n480_), .C2(new_n472_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n482_), .A2(new_n484_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT70), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n484_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT73), .ZN(new_n497_));
  INV_X1    g296(.A(G22gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n347_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G15gat), .A2(G22gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G1gat), .A2(G8gat), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n499_), .A2(new_n500_), .B1(KEYINPUT14), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n497_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT74), .Z(new_n510_));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n503_), .B(new_n507_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n510_), .A2(new_n513_), .B1(new_n514_), .B2(new_n512_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G113gat), .B(G141gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT75), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G169gat), .B(G197gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n495_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n434_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n462_), .A2(new_n507_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n508_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n525_), .B(new_n526_), .C1(KEYINPUT35), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n531_), .A2(KEYINPUT36), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(KEYINPUT36), .Z(new_n536_));
  AND2_X1   g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n536_), .B(KEYINPUT71), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n531_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT37), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n463_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n503_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT16), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n547_), .A2(new_n553_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n544_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n524_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G1gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n411_), .B(KEYINPUT98), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT38), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(KEYINPUT100), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(KEYINPUT38), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(KEYINPUT100), .A3(new_n565_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n538_), .A2(new_n558_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n524_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n411_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G1gat), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n573_), .A2(KEYINPUT99), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(KEYINPUT99), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n568_), .B(new_n569_), .C1(new_n574_), .C2(new_n575_), .ZN(G1324gat));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n319_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n337_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n335_), .A2(KEYINPUT96), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n325_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT97), .B1(new_n581_), .B2(new_n324_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n342_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n524_), .A2(new_n584_), .A3(new_n570_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT101), .B1(new_n585_), .B2(G8gat), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT102), .B(new_n577_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G8gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n560_), .A2(new_n593_), .A3(new_n584_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n589_), .A2(new_n592_), .A3(KEYINPUT40), .A4(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1325gat));
  NAND3_X1  g398(.A1(new_n560_), .A2(new_n347_), .A3(new_n413_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n571_), .A2(new_n413_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n601_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT41), .B1(new_n601_), .B2(G15gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(G1326gat));
  NAND3_X1  g403(.A1(new_n560_), .A2(new_n498_), .A3(new_n250_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n571_), .A2(new_n250_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G22gat), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(G1327gat));
  NOR3_X1   g409(.A1(new_n535_), .A2(new_n537_), .A3(new_n557_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n524_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n411_), .ZN(new_n613_));
  OR3_X1    g412(.A1(new_n612_), .A2(G29gat), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n523_), .A2(new_n557_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n249_), .B(new_n412_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n416_), .A2(new_n420_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT94), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(new_n249_), .A3(new_n431_), .A4(new_n428_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n433_), .A2(new_n373_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n616_), .B1(new_n622_), .B2(new_n544_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n540_), .A2(new_n543_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT43), .B(new_n624_), .C1(new_n617_), .C2(new_n621_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n615_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n434_), .B2(new_n624_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n616_), .A3(new_n544_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(KEYINPUT44), .A3(new_n615_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n563_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT103), .B1(new_n634_), .B2(G29gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n614_), .B1(new_n635_), .B2(new_n636_), .ZN(G1328gat));
  AND2_X1   g436(.A1(new_n584_), .A2(KEYINPUT104), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n584_), .A2(KEYINPUT104), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n612_), .A2(G36gat), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n628_), .A2(new_n584_), .A3(new_n632_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G36gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT46), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n645_), .A3(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1329gat));
  INV_X1    g449(.A(G43gat), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n373_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n628_), .A2(new_n632_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n628_), .A2(new_n632_), .A3(KEYINPUT105), .A4(new_n652_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n612_), .B2(new_n373_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .A4(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1330gat));
  INV_X1    g462(.A(new_n612_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G50gat), .B1(new_n664_), .B2(new_n250_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n250_), .A2(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n633_), .B2(new_n666_), .ZN(G1331gat));
  AOI211_X1 g466(.A(new_n522_), .B(new_n495_), .C1(new_n617_), .C2(new_n621_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n559_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT107), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT107), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n563_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n522_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n557_), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n434_), .A2(new_n495_), .A3(new_n538_), .A4(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n613_), .A2(new_n673_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n672_), .A2(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1332gat));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n640_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n640_), .A2(G64gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT109), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n669_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n676_), .B2(new_n413_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NOR2_X1   g488(.A1(new_n373_), .A2(G71gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT110), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n669_), .B2(new_n691_), .ZN(G1334gat));
  AOI21_X1  g491(.A(new_n229_), .B1(new_n676_), .B2(new_n250_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT50), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n250_), .A2(new_n229_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT111), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n669_), .B2(new_n696_), .ZN(G1335gat));
  NAND2_X1  g496(.A1(new_n668_), .A2(new_n611_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n668_), .A2(KEYINPUT112), .A3(new_n611_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G85gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n563_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n631_), .A2(KEYINPUT113), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n629_), .A2(new_n706_), .A3(new_n630_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT114), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n522_), .A2(new_n557_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n489_), .A2(new_n494_), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n489_), .A2(new_n494_), .A3(new_n709_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT114), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n705_), .A2(new_n707_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n411_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n704_), .B1(new_n714_), .B2(new_n703_), .ZN(G1336gat));
  INV_X1    g514(.A(G92gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n702_), .A2(new_n716_), .A3(new_n584_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n713_), .A2(new_n680_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n716_), .ZN(G1337gat));
  AOI21_X1  g518(.A(new_n450_), .B1(new_n713_), .B2(new_n413_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n702_), .A2(new_n413_), .A3(new_n442_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(KEYINPUT115), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n702_), .A2(new_n231_), .A3(new_n250_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n712_), .A2(new_n710_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n250_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G106gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n249_), .B1(new_n712_), .B2(new_n710_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT116), .A3(new_n733_), .A4(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n733_), .B1(new_n737_), .B2(G106gat), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n735_), .B(new_n738_), .C1(new_n739_), .C2(KEYINPUT117), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT117), .B(KEYINPUT52), .C1(new_n732_), .C2(new_n231_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n727_), .B(new_n728_), .C1(new_n740_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n732_), .B2(new_n231_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n747_), .A2(new_n741_), .A3(new_n735_), .A4(new_n738_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n728_), .B1(new_n748_), .B2(new_n727_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n744_), .A2(new_n749_), .ZN(G1339gat));
  INV_X1    g549(.A(G113gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n461_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT55), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n480_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT55), .B(new_n469_), .C1(new_n461_), .C2(new_n465_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n471_), .A2(new_n754_), .A3(KEYINPUT55), .ZN(new_n759_));
  INV_X1    g558(.A(new_n757_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT119), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n478_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT120), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n752_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n479_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n674_), .A2(new_n765_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n756_), .A2(new_n753_), .A3(new_n757_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT119), .B1(new_n759_), .B2(new_n760_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n477_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n764_), .B(new_n766_), .C1(new_n770_), .C2(new_n763_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n511_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n510_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n519_), .B1(new_n514_), .B2(new_n511_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n521_), .A2(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n490_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n538_), .B1(new_n771_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n762_), .A2(new_n752_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n776_), .A2(new_n765_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n770_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n544_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n781_), .A2(new_n782_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n778_), .A2(KEYINPUT57), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n787_), .B(new_n538_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n558_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n544_), .A2(new_n675_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT54), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n373_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n343_), .A2(new_n563_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n751_), .B1(new_n795_), .B2(new_n674_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT121), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n751_), .C1(new_n795_), .C2(new_n674_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n793_), .A2(KEYINPUT59), .A3(new_n794_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n674_), .A2(new_n751_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n797_), .A2(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(G1340gat));
  INV_X1    g604(.A(new_n795_), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n495_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n806_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n807_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n495_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n807_), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n795_), .B2(new_n558_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT122), .B(new_n812_), .C1(new_n795_), .C2(new_n558_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n558_), .A2(new_n812_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n815_), .A2(new_n816_), .B1(new_n803_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g617(.A(G134gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n806_), .A2(new_n819_), .A3(new_n538_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n624_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(G1343gat));
  NOR2_X1   g621(.A1(new_n413_), .A2(new_n249_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n680_), .A2(new_n562_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n522_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G141gat), .ZN(G1344gat));
  AND2_X1   g628(.A1(new_n489_), .A2(new_n494_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g631(.A1(new_n789_), .A2(new_n792_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(new_n557_), .A3(new_n823_), .A4(new_n826_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT123), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n825_), .A2(new_n836_), .A3(new_n557_), .A4(new_n826_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n835_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(G162gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n827_), .A2(new_n842_), .A3(new_n538_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n827_), .A2(new_n544_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1347gat));
  NOR3_X1   g644(.A1(new_n640_), .A2(new_n250_), .A3(new_n563_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n833_), .A2(new_n413_), .A3(new_n522_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G169gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n793_), .A2(new_n297_), .A3(new_n522_), .A4(new_n846_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n849_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(G1348gat));
  NAND2_X1  g652(.A1(new_n793_), .A2(new_n846_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n495_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n268_), .ZN(G1349gat));
  NAND3_X1  g655(.A1(new_n793_), .A2(new_n557_), .A3(new_n846_), .ZN(new_n857_));
  MUX2_X1   g656(.A(new_n280_), .B(G183gat), .S(new_n857_), .Z(G1350gat));
  INV_X1    g657(.A(KEYINPUT125), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n833_), .A2(new_n413_), .A3(new_n544_), .A4(new_n846_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n860_), .A2(G190gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n538_), .A2(new_n281_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n854_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n859_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(G190gat), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(KEYINPUT125), .C1(new_n854_), .C2(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1351gat));
  NOR2_X1   g666(.A1(new_n640_), .A2(new_n411_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n825_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n522_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n830_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G204gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT126), .B(G204gat), .Z(new_n875_));
  NAND3_X1  g674(.A1(new_n869_), .A2(new_n830_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1353gat));
  NOR3_X1   g676(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n558_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n869_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n880_), .B(new_n882_), .ZN(G1354gat));
  INV_X1    g682(.A(G218gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n869_), .A2(new_n884_), .A3(new_n538_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n869_), .A2(new_n544_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1355gat));
endmodule


