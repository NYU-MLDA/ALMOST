//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT86), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT2), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n211_), .B(new_n212_), .C1(new_n213_), .C2(new_n205_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n203_), .B(new_n204_), .C1(new_n208_), .C2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n203_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n207_), .A2(new_n209_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  OR3_X1    g020(.A1(new_n221_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G22gat), .B(G50gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT89), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G228gat), .A2(G233gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(G197gat), .B(G204gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT87), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n228_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n215_), .A2(new_n220_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n236_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n241_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G78gat), .B(G106gat), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n227_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n227_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n225_), .A2(new_n226_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n245_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(KEYINPUT90), .ZN(new_n256_));
  OAI22_X1  g055(.A1(new_n249_), .A2(new_n251_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT23), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  INV_X1    g060(.A(G169gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT22), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(KEYINPUT22), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n263_), .A2(new_n264_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n260_), .B(new_n261_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT25), .B(G183gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT81), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n275_), .B(new_n259_), .C1(KEYINPUT24), .C2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n270_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G71gat), .B(G99gat), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n284_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT84), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n288_), .B(new_n289_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT84), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT30), .B(G15gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT31), .B(G43gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n287_), .B(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n257_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n240_), .A2(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n221_), .A2(new_n292_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT4), .B1(new_n221_), .B2(new_n292_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n301_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT4), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(new_n305_), .B2(new_n300_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307_));
  INV_X1    g106(.A(G85gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n302_), .B(new_n313_), .C1(new_n305_), .C2(new_n300_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT95), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n236_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n276_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n259_), .B1(KEYINPUT24), .B2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT91), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(KEYINPUT91), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n328_), .A2(new_n279_), .A3(new_n273_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n263_), .A2(new_n267_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n260_), .B(new_n261_), .C1(G176gat), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n325_), .B1(new_n335_), .B2(new_n236_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n236_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n334_), .A3(new_n330_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n282_), .A2(new_n236_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT20), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n338_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n324_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n282_), .A2(new_n236_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n334_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n330_), .A2(new_n331_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n331_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(KEYINPUT20), .B(new_n347_), .C1(new_n351_), .C2(new_n341_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n341_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n339_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n352_), .A2(new_n338_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n346_), .A2(KEYINPUT96), .B1(new_n322_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n352_), .A2(new_n338_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n345_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n323_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT96), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n317_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n322_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n336_), .A2(new_n339_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n353_), .A2(new_n354_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n355_), .A2(new_n322_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n317_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n298_), .B(new_n316_), .C1(new_n362_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT97), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n257_), .A2(new_n297_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT96), .B(new_n323_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n367_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n346_), .A2(KEYINPUT96), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT27), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT97), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n316_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  INV_X1    g179(.A(new_n300_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n305_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n299_), .A2(new_n381_), .A3(new_n301_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n382_), .A2(new_n311_), .A3(new_n383_), .ZN(new_n384_));
  OR3_X1    g183(.A1(new_n305_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n314_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n314_), .A2(new_n387_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n366_), .A2(new_n367_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n364_), .A2(new_n365_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n395_), .A2(new_n316_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n257_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n361_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n369_), .B1(new_n399_), .B2(KEYINPUT27), .ZN(new_n400_));
  OAI221_X1 g199(.A(new_n316_), .B1(new_n253_), .B2(new_n256_), .C1(new_n249_), .C2(new_n251_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n297_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n371_), .A2(new_n379_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G43gat), .B(G50gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT74), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G15gat), .B(G22gat), .ZN(new_n409_));
  INV_X1    g208(.A(G1gat), .ZN(new_n410_));
  INV_X1    g209(.A(G8gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT14), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G8gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n408_), .B(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n408_), .A2(new_n416_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G229gat), .A2(G233gat), .ZN(new_n421_));
  MUX2_X1   g220(.A(new_n417_), .B(new_n420_), .S(new_n421_), .Z(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n422_), .A2(KEYINPUT79), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n422_), .B2(KEYINPUT79), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G57gat), .B(G64gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT69), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n434_));
  XOR2_X1   g233(.A(G71gat), .B(G78gat), .Z(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n432_), .A2(KEYINPUT69), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(KEYINPUT69), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n438_), .A2(new_n439_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT12), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n445_));
  INV_X1    g244(.A(G99gat), .ZN(new_n446_));
  INV_X1    g245(.A(G106gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n444_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT8), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT8), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459_));
  AND3_X1   g258(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n453_), .A2(KEYINPUT65), .A3(new_n454_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n450_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n458_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI211_X1 g265(.A(KEYINPUT67), .B(new_n450_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n457_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT64), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n446_), .A2(KEYINPUT10), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT10), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G99gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n473_), .B2(new_n447_), .ZN(new_n474_));
  AOI211_X1 g273(.A(KEYINPUT64), .B(G106gat), .C1(new_n470_), .C2(new_n472_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n462_), .A2(new_n463_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n444_), .B2(KEYINPUT9), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT66), .B1(new_n476_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT10), .B(G99gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT64), .B1(new_n483_), .B2(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n469_), .A3(new_n447_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n441_), .B1(new_n468_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n468_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT68), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n468_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n437_), .A2(new_n440_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n496_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n489_), .A2(new_n493_), .A3(new_n468_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n493_), .B1(new_n489_), .B2(new_n468_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n496_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n500_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G120gat), .B(G148gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G176gat), .B(G204gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT71), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n503_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT72), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n520_), .A2(new_n522_), .A3(KEYINPUT13), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT13), .B1(new_n520_), .B2(new_n522_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n404_), .A2(new_n430_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n495_), .A2(new_n408_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n419_), .B2(new_n491_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT75), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT73), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n527_), .A2(new_n531_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n532_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT37), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n543_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT76), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n415_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(new_n496_), .Z(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT17), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT16), .B(G183gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  MUX2_X1   g360(.A(KEYINPUT17), .B(new_n557_), .S(new_n561_), .Z(new_n562_));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n556_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n552_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT78), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n526_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n410_), .A3(new_n315_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n549_), .A2(new_n543_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n568_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n526_), .A2(new_n315_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(G1gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n582_), .ZN(G1324gat));
  NAND3_X1  g382(.A1(new_n526_), .A2(new_n400_), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(G8gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT39), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n411_), .A3(new_n400_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n588_), .B(new_n590_), .ZN(G1325gat));
  OR3_X1    g390(.A1(new_n572_), .A2(G15gat), .A3(new_n403_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n526_), .A2(new_n297_), .A3(new_n580_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n593_), .A2(G15gat), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n593_), .B2(G15gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT101), .ZN(G1326gat));
  OR3_X1    g397(.A1(new_n572_), .A2(G22gat), .A3(new_n257_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n257_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n526_), .A2(new_n600_), .A3(new_n580_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G22gat), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT42), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT42), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n599_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT102), .Z(G1327gat));
  NOR2_X1   g405(.A1(new_n569_), .A2(new_n578_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n526_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(G29gat), .B1(new_n608_), .B2(new_n315_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT43), .B1(new_n404_), .B2(new_n552_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n401_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n397_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n384_), .A2(new_n385_), .B1(new_n387_), .B2(new_n314_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n613_), .A2(new_n367_), .A3(new_n366_), .A4(new_n388_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n600_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n403_), .B1(new_n611_), .B2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n370_), .A2(KEYINPUT97), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n378_), .B1(new_n377_), .B2(new_n316_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  INV_X1    g419(.A(new_n552_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n569_), .B1(new_n610_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT44), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n525_), .A2(new_n430_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(KEYINPUT44), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n628_), .A3(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n315_), .A2(G29gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n609_), .B1(new_n632_), .B2(new_n633_), .ZN(G1328gat));
  INV_X1    g433(.A(G36gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n400_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT104), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT104), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n608_), .A2(new_n635_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT45), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n635_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n641_), .B(KEYINPUT46), .C1(new_n635_), .C2(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  INV_X1    g446(.A(KEYINPUT47), .ZN(new_n648_));
  INV_X1    g447(.A(new_n631_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n628_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n297_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G43gat), .ZN(new_n652_));
  INV_X1    g451(.A(G43gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n608_), .A2(new_n653_), .A3(new_n297_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n648_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n403_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n648_), .B(new_n654_), .C1(new_n656_), .C2(new_n653_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1330gat));
  INV_X1    g458(.A(G50gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n608_), .A2(new_n660_), .A3(new_n600_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n257_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT105), .ZN(new_n663_));
  OAI21_X1  g462(.A(G50gat), .B1(new_n662_), .B2(KEYINPUT105), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(G1331gat));
  NAND2_X1  g464(.A1(new_n525_), .A2(new_n430_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n404_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n580_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(G57gat), .A3(new_n315_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n571_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G57gat), .B1(new_n673_), .B2(new_n315_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(G1332gat));
  INV_X1    g474(.A(G64gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n668_), .B2(new_n639_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT48), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n639_), .A2(new_n676_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT107), .Z(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n672_), .B2(new_n680_), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n668_), .B2(new_n297_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT49), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n682_), .A3(new_n297_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n668_), .B2(new_n600_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT50), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n673_), .A2(new_n687_), .A3(new_n600_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1335gat));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n610_), .A2(new_n622_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n666_), .A2(new_n569_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n610_), .B2(new_n622_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n610_), .A2(new_n622_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT108), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n315_), .A2(G85gat), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT110), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n667_), .A2(new_n607_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n308_), .B1(new_n705_), .B2(new_n316_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1336gat));
  AND4_X1   g508(.A1(G92gat), .A2(new_n697_), .A3(new_n639_), .A4(new_n701_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n705_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G92gat), .B1(new_n711_), .B2(new_n400_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1337gat));
  NAND3_X1  g512(.A1(new_n697_), .A2(new_n297_), .A3(new_n701_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G99gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(new_n473_), .A3(new_n297_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n719_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1338gat));
  NOR3_X1   g520(.A1(new_n705_), .A2(G106gat), .A3(new_n257_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT112), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n623_), .A2(new_n430_), .A3(new_n525_), .A4(new_n600_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(new_n725_), .A3(G106gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G106gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g528(.A1(new_n429_), .A2(new_n518_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT56), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n498_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT113), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n504_), .A2(new_n505_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT12), .B1(new_n735_), .B2(new_n499_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n499_), .A2(KEYINPUT12), .A3(new_n491_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n506_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n508_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(KEYINPUT55), .ZN(new_n741_));
  INV_X1    g540(.A(new_n503_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n734_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n516_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n734_), .B2(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n731_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n734_), .A2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n503_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n516_), .A4(new_n743_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n730_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  MUX2_X1   g549(.A(new_n420_), .B(new_n417_), .S(new_n421_), .Z(new_n751_));
  MUX2_X1   g550(.A(new_n422_), .B(new_n751_), .S(new_n425_), .Z(new_n752_));
  AND3_X1   g551(.A1(new_n520_), .A2(new_n522_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n578_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(KEYINPUT114), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n746_), .A2(new_n749_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n518_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n760_), .A2(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n764_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n761_), .C1(new_n746_), .C2(new_n749_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n621_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT57), .B(new_n578_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n758_), .A2(new_n759_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n568_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n525_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n429_), .B(new_n568_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n771_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n400_), .A2(new_n316_), .A3(new_n372_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G113gat), .B1(new_n783_), .B2(new_n429_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n768_), .A2(new_n756_), .A3(new_n769_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n568_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n778_), .B1(new_n786_), .B2(KEYINPUT116), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(new_n568_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n400_), .A2(KEYINPUT59), .A3(new_n316_), .A4(new_n372_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n782_), .A2(KEYINPUT59), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(G113gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n429_), .A2(KEYINPUT117), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G113gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n784_), .B1(new_n792_), .B2(new_n796_), .ZN(G1340gat));
  AND2_X1   g596(.A1(new_n792_), .A2(new_n525_), .ZN(new_n798_));
  INV_X1    g597(.A(G120gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n800_));
  AOI21_X1  g599(.A(G120gat), .B1(new_n525_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n801_), .A2(new_n802_), .B1(KEYINPUT60), .B2(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n802_), .B2(new_n801_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n783_), .A2(KEYINPUT119), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT119), .B1(new_n783_), .B2(new_n804_), .ZN(new_n806_));
  OAI22_X1  g605(.A1(new_n798_), .A2(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(G1341gat));
  AOI21_X1  g606(.A(G127gat), .B1(new_n783_), .B2(new_n569_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n569_), .A2(G127gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n792_), .B2(new_n809_), .ZN(G1342gat));
  AOI21_X1  g609(.A(G134gat), .B1(new_n783_), .B2(new_n579_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n621_), .A2(G134gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n792_), .B2(new_n812_), .ZN(G1343gat));
  AOI21_X1  g612(.A(new_n778_), .B1(new_n770_), .B2(new_n568_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n257_), .A2(new_n297_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR4_X1   g615(.A1(new_n814_), .A2(new_n316_), .A3(new_n639_), .A4(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n429_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT120), .B(G141gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1344gat));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n525_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n569_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  AOI21_X1  g624(.A(G162gat), .B1(new_n817_), .B2(new_n579_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n621_), .A2(G162gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n817_), .B2(new_n827_), .ZN(G1347gat));
  NAND2_X1  g627(.A1(new_n639_), .A2(new_n316_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n372_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n430_), .B(new_n831_), .C1(new_n787_), .C2(new_n789_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT121), .B(KEYINPUT62), .C1(new_n832_), .C2(new_n262_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n790_), .A2(new_n429_), .A3(new_n830_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(G169gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(G169gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT121), .B1(new_n839_), .B2(KEYINPUT62), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n833_), .B1(new_n838_), .B2(new_n840_), .ZN(G1348gat));
  NAND2_X1  g640(.A1(new_n790_), .A2(new_n830_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n266_), .B1(new_n842_), .B2(new_n772_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n780_), .A2(KEYINPUT122), .A3(new_n257_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n814_), .B2(new_n600_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n829_), .A2(new_n403_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n772_), .A2(new_n266_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .A4(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n843_), .A2(new_n849_), .A3(KEYINPUT123), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1349gat));
  NOR3_X1   g653(.A1(new_n842_), .A2(new_n271_), .A3(new_n568_), .ZN(new_n855_));
  INV_X1    g654(.A(G183gat), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n844_), .A2(new_n846_), .A3(new_n569_), .A4(new_n847_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n842_), .B2(new_n552_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n579_), .A2(new_n272_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n842_), .B2(new_n860_), .ZN(G1351gat));
  NOR3_X1   g660(.A1(new_n814_), .A2(new_n816_), .A3(new_n829_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n862_), .A2(new_n429_), .B1(KEYINPUT124), .B2(G197gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n863_), .B(new_n864_), .Z(G1352gat));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n525_), .ZN(new_n866_));
  INV_X1    g665(.A(G204gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(KEYINPUT125), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n867_), .A2(KEYINPUT125), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n866_), .B2(new_n868_), .ZN(G1353gat));
  INV_X1    g670(.A(KEYINPUT63), .ZN(new_n872_));
  INV_X1    g671(.A(new_n829_), .ZN(new_n873_));
  INV_X1    g672(.A(G211gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n569_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT126), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n780_), .A2(new_n815_), .A3(new_n873_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n814_), .A2(new_n816_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n873_), .A4(new_n876_), .ZN(new_n881_));
  AND4_X1   g680(.A1(new_n872_), .A2(new_n878_), .A3(new_n874_), .A4(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n878_), .A2(new_n881_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1354gat));
  AOI21_X1  g683(.A(G218gat), .B1(new_n862_), .B2(new_n579_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n621_), .A2(G218gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n862_), .B2(new_n886_), .ZN(G1355gat));
endmodule


