//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT92), .Z(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT96), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT3), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT93), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n209_), .C1(KEYINPUT2), .C2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(KEYINPUT95), .A3(KEYINPUT1), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT95), .B1(new_n213_), .B2(KEYINPUT1), .ZN(new_n217_));
  OAI221_X1 g016(.A(new_n214_), .B1(KEYINPUT1), .B2(new_n213_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n208_), .B(KEYINPUT94), .Z(new_n219_));
  INV_X1    g018(.A(new_n211_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT4), .B1(new_n205_), .B2(new_n222_), .ZN(new_n223_));
  MUX2_X1   g022(.A(new_n204_), .B(new_n205_), .S(new_n222_), .Z(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(KEYINPUT4), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT33), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G1gat), .B(G29gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G85gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G57gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  NAND4_X1  g033(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .A4(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n230_), .B(new_n234_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT33), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G8gat), .B(G36gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT18), .B(G64gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(G190gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT23), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT89), .ZN(new_n248_));
  OR3_X1    g047(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT23), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(KEYINPUT25), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n245_), .A2(KEYINPUT25), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n256_), .A2(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n252_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n249_), .A2(new_n247_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n245_), .A2(new_n246_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265_));
  AOI21_X1  g064(.A(G176gat), .B1(new_n265_), .B2(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT22), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n263_), .A2(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT86), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n260_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT100), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(KEYINPUT100), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n262_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT97), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT21), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G197gat), .B(G204gat), .Z(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n279_), .C1(KEYINPUT21), .C2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n250_), .A2(new_n264_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n265_), .A2(KEYINPUT87), .A3(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n268_), .A2(KEYINPUT87), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n266_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n271_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n255_), .B(KEYINPUT85), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n253_), .B(KEYINPUT84), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n257_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n251_), .B1(new_n271_), .B2(new_n259_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n263_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n282_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n286_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n293_), .A2(new_n298_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n275_), .A2(new_n282_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT20), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n285_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT101), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT101), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n304_), .B2(new_n285_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n244_), .B(new_n301_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(KEYINPUT101), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n301_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n243_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n224_), .A2(new_n226_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n234_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n313_), .B(new_n314_), .C1(new_n225_), .C2(new_n229_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n238_), .A2(new_n309_), .A3(new_n312_), .A4(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n230_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n236_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n244_), .A2(KEYINPUT32), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n283_), .A2(KEYINPUT102), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n283_), .A2(KEYINPUT102), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n300_), .A3(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n323_), .A2(KEYINPUT103), .A3(new_n285_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n285_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n302_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n303_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n323_), .A2(new_n285_), .B1(KEYINPUT103), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n320_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n319_), .B(new_n328_), .C1(new_n311_), .C2(new_n320_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n316_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT31), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n205_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(new_n299_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G15gat), .B(G43gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n337_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n334_), .B(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G78gat), .B(G106gat), .Z(new_n342_));
  OR3_X1    g141(.A1(new_n222_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n282_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n282_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n349_), .B(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n342_), .B1(new_n347_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT99), .B1(new_n347_), .B2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n346_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n345_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n353_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n342_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n330_), .A2(new_n341_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n319_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n341_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n334_), .B(new_n340_), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n354_), .A2(new_n360_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT99), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n372_), .B2(new_n361_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n366_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n243_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT104), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n310_), .A2(new_n376_), .A3(new_n244_), .A4(new_n301_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n309_), .A2(KEYINPUT104), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT27), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT27), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n312_), .A2(new_n381_), .A3(new_n309_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n365_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT76), .B(G15gat), .ZN(new_n387_));
  INV_X1    g186(.A(G22gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G1gat), .ZN(new_n390_));
  INV_X1    g189(.A(G8gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT14), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G8gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT77), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n395_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G43gat), .B(G50gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(G29gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G229gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT15), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n401_), .B(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n398_), .B(new_n401_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n411_), .B2(new_n404_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n412_), .B2(new_n408_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n386_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT81), .B(G113gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G141gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G169gat), .B(G197gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT80), .B1(new_n420_), .B2(KEYINPUT83), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n415_), .A2(new_n420_), .B1(new_n421_), .B2(new_n413_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n385_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT105), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT11), .ZN(new_n427_));
  INV_X1    g226(.A(G78gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G71gat), .ZN(new_n429_));
  INV_X1    g228(.A(G71gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G78gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G57gat), .A2(G64gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G57gat), .A2(G64gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT68), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G57gat), .ZN(new_n436_));
  INV_X1    g235(.A(G64gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G57gat), .A2(G64gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI211_X1 g240(.A(new_n427_), .B(new_n432_), .C1(new_n435_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n427_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n435_), .A2(new_n441_), .A3(new_n427_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n432_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G85gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n240_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n451_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT65), .A3(G85gat), .A4(G92gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT10), .B(G99gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT64), .B(G106gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n460_), .B(new_n463_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n450_), .A2(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n461_), .A2(KEYINPUT8), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n451_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n457_), .A2(new_n459_), .A3(KEYINPUT66), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT66), .B1(new_n457_), .B2(new_n459_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT67), .A3(new_n452_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n475_), .B1(new_n478_), .B2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n443_), .B(new_n447_), .C1(new_n472_), .C2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n458_), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n457_), .A2(new_n459_), .A3(KEYINPUT66), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n484_), .A2(KEYINPUT67), .A3(new_n452_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n452_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n495_), .B(new_n496_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n474_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n451_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n460_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n484_), .A2(new_n452_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n473_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n466_), .A2(new_n471_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n435_), .A2(new_n441_), .A3(new_n427_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n444_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n442_), .B1(new_n509_), .B2(new_n432_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n491_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n472_), .A2(new_n487_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n447_), .A2(new_n443_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT69), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(KEYINPUT70), .A3(new_n510_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n490_), .A2(new_n511_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT71), .B1(new_n512_), .B2(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT12), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n513_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n488_), .A2(KEYINPUT71), .A3(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n521_), .A2(new_n517_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n519_), .B2(new_n525_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n519_), .A2(new_n525_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n530_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n532_), .A3(new_n531_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n539_), .A3(KEYINPUT13), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n385_), .A2(KEYINPUT105), .A3(new_n423_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n426_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n507_), .A2(new_n401_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n406_), .B2(new_n507_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT35), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT75), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(KEYINPUT35), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n552_), .B(KEYINPUT75), .C1(new_n554_), .C2(new_n548_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G218gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT74), .B(G190gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n553_), .A2(new_n555_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n564_), .A2(KEYINPUT37), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT37), .B1(new_n564_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n398_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n513_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT16), .B(G183gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n572_), .A2(KEYINPUT78), .A3(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n572_), .A2(new_n580_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n571_), .A2(new_n510_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n571_), .A2(new_n510_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n577_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n569_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n546_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n390_), .A3(new_n319_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n564_), .A2(new_n565_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n588_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n383_), .B(new_n366_), .C1(new_n373_), .C2(new_n367_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n365_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n544_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n422_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n366_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n602_), .ZN(G1324gat));
  XNOR2_X1  g402(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT110), .ZN(new_n606_));
  INV_X1    g405(.A(new_n596_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n385_), .A2(new_n600_), .A3(new_n384_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT107), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT108), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT107), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n598_), .A2(new_n612_), .A3(new_n600_), .A4(new_n384_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n609_), .A2(G8gat), .A3(new_n611_), .A4(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(KEYINPUT108), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n546_), .A2(new_n391_), .A3(new_n384_), .A4(new_n590_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n606_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n609_), .A2(new_n613_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(G8gat), .A3(new_n615_), .A4(new_n611_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(KEYINPUT108), .A3(new_n610_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n606_), .A2(new_n620_), .A3(new_n617_), .A4(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n605_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n606_), .A3(new_n617_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT110), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n626_), .A3(new_n604_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n601_), .B2(new_n341_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT41), .Z(new_n630_));
  INV_X1    g429(.A(new_n591_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n341_), .A2(G15gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n601_), .B2(new_n364_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(new_n364_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n388_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n631_), .B2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n595_), .A2(new_n588_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n426_), .A2(new_n544_), .A3(new_n545_), .A4(new_n639_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n640_), .A2(G29gat), .A3(new_n366_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n385_), .A2(new_n569_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT43), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n385_), .A2(new_n644_), .A3(new_n569_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n600_), .A3(new_n589_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n646_), .A2(KEYINPUT44), .A3(new_n600_), .A4(new_n589_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n319_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT111), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n651_), .A2(new_n652_), .A3(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n651_), .B2(G29gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n641_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n384_), .A3(new_n650_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(G36gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n640_), .A2(G36gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n384_), .ZN(new_n661_));
  NOR4_X1   g460(.A1(new_n640_), .A2(KEYINPUT45), .A3(G36gat), .A4(new_n383_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(G36gat), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(KEYINPUT46), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1329gat));
  NAND4_X1  g466(.A1(new_n649_), .A2(G43gat), .A3(new_n368_), .A4(new_n650_), .ZN(new_n668_));
  INV_X1    g467(.A(G43gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n640_), .B2(new_n341_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g471(.A1(new_n649_), .A2(new_n636_), .A3(new_n650_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G50gat), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n640_), .A2(G50gat), .A3(new_n364_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT112), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT112), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n544_), .A2(new_n423_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n385_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n590_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT113), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n319_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n682_), .A2(new_n607_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n319_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(G57gat), .B2(new_n687_), .ZN(G1332gat));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n437_), .A3(new_n384_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n686_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G64gat), .B1(new_n690_), .B2(new_n383_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT48), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT48), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT114), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT114), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n689_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1333gat));
  AOI21_X1  g497(.A(new_n430_), .B1(new_n686_), .B2(new_n368_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT49), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n684_), .A2(new_n430_), .A3(new_n368_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1334gat));
  AOI21_X1  g501(.A(new_n428_), .B1(new_n686_), .B2(new_n636_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT50), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n684_), .A2(new_n428_), .A3(new_n636_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  AND2_X1   g505(.A1(new_n682_), .A2(new_n639_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n319_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT115), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n646_), .A2(new_n589_), .A3(new_n681_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n366_), .A2(new_n448_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  AOI21_X1  g511(.A(G92gat), .B1(new_n707_), .B2(new_n384_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n710_), .A2(G92gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n384_), .ZN(G1337gat));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n368_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n341_), .A2(new_n464_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n716_), .A2(G99gat), .B1(new_n707_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(G1338gat));
  INV_X1    g519(.A(new_n465_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n707_), .A2(new_n721_), .A3(new_n636_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n646_), .A2(new_n636_), .A3(new_n589_), .A4(new_n681_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1339gat));
  NOR2_X1   g528(.A1(new_n384_), .A2(new_n366_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT57), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n413_), .A2(new_n420_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n411_), .A2(new_n404_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n403_), .A2(new_n407_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(G229gat), .A3(G233gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n420_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n540_), .A2(new_n733_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT120), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n518_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(KEYINPUT55), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT119), .B(new_n744_), .C1(new_n741_), .C2(new_n518_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n525_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT71), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n747_), .B(KEYINPUT12), .C1(new_n507_), .C2(new_n510_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n523_), .B1(new_n488_), .B2(KEYINPUT71), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n517_), .B1(new_n750_), .B2(new_n522_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT119), .B1(new_n751_), .B2(new_n744_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n525_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n740_), .A3(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n755_), .A3(new_n537_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n739_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n746_), .A2(new_n755_), .A3(KEYINPUT56), .A4(new_n537_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n422_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n756_), .A2(KEYINPUT120), .A3(new_n757_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n531_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n738_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n595_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n732_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n756_), .A2(new_n757_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT120), .A3(new_n759_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n746_), .A2(new_n755_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(new_n739_), .A3(KEYINPUT56), .A4(new_n537_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n768_), .A2(new_n423_), .A3(new_n531_), .A4(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n738_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT57), .A3(new_n595_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n767_), .A2(new_n759_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n733_), .A2(new_n737_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n531_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n775_), .A2(KEYINPUT58), .A3(new_n531_), .A4(new_n776_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n569_), .A3(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n766_), .A2(new_n774_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n589_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n543_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT13), .B1(new_n535_), .B2(new_n539_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n422_), .B(new_n588_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n544_), .A2(KEYINPUT117), .A3(new_n422_), .A4(new_n588_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n790_), .A2(new_n568_), .A3(new_n793_), .A4(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n789_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n791_), .B(new_n792_), .C1(new_n796_), .C2(new_n569_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n731_), .B1(new_n783_), .B2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n367_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n423_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n803_), .A3(new_n367_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n800_), .B2(new_n367_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n802_), .B1(new_n807_), .B2(new_n423_), .ZN(G1340gat));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT121), .B1(new_n809_), .B2(KEYINPUT60), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n801_), .B(new_n812_), .C1(new_n813_), .C2(new_n810_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n804_), .A2(new_n805_), .A3(new_n544_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n801_), .B2(new_n588_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n804_), .A2(new_n805_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n588_), .A2(G127gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(G1342gat));
  AOI21_X1  g619(.A(G134gat), .B1(new_n801_), .B2(new_n765_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n569_), .A2(G134gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n818_), .B2(new_n822_), .ZN(G1343gat));
  NAND2_X1  g622(.A1(new_n783_), .A2(new_n799_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n373_), .A3(new_n730_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT122), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n800_), .A2(new_n827_), .A3(new_n373_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G141gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n423_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n827_), .B1(new_n800_), .B2(new_n373_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n798_), .B1(new_n782_), .B2(new_n589_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n373_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n833_), .A2(KEYINPUT122), .A3(new_n834_), .A4(new_n731_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n423_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G141gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n837_), .ZN(G1344gat));
  XNOR2_X1  g637(.A(KEYINPUT123), .B(G148gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n829_), .B2(new_n599_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n599_), .B(new_n839_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1345gat));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n829_), .B2(new_n588_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n588_), .B(new_n844_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1346gat));
  AOI21_X1  g647(.A(G162gat), .B1(new_n829_), .B2(new_n765_), .ZN(new_n849_));
  OAI211_X1 g648(.A(G162gat), .B(new_n569_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1347gat));
  XOR2_X1   g651(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n833_), .A2(new_n319_), .A3(new_n383_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n855_), .A2(new_n423_), .A3(new_n367_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n267_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n265_), .A2(G169gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n858_), .A3(new_n268_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n367_), .ZN(new_n860_));
  OAI211_X1 g659(.A(G169gat), .B(new_n853_), .C1(new_n860_), .C2(new_n422_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n859_), .A3(new_n861_), .ZN(G1348gat));
  NAND3_X1  g661(.A1(new_n855_), .A2(new_n599_), .A3(new_n367_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g663(.A1(new_n860_), .A2(new_n256_), .A3(new_n589_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n588_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n245_), .B2(new_n867_), .ZN(G1350gat));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n257_), .A3(new_n765_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G190gat), .B1(new_n860_), .B2(new_n568_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1351gat));
  NAND3_X1  g670(.A1(new_n855_), .A2(new_n423_), .A3(new_n373_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT125), .B(G197gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1352gat));
  NAND3_X1  g673(.A1(new_n855_), .A2(new_n599_), .A3(new_n373_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT127), .Z(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n589_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT126), .Z(new_n881_));
  NAND3_X1  g680(.A1(new_n855_), .A2(new_n373_), .A3(new_n881_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n878_), .B(new_n879_), .S(new_n882_), .Z(G1354gat));
  AND3_X1   g682(.A1(new_n855_), .A2(new_n373_), .A3(new_n765_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n855_), .A2(new_n373_), .A3(new_n569_), .ZN(new_n885_));
  MUX2_X1   g684(.A(new_n884_), .B(new_n885_), .S(G218gat), .Z(G1355gat));
endmodule


