//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(G233gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT91), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT91), .ZN(new_n204_));
  OAI21_X1  g003(.A(G228gat), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206_));
  AND2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n214_));
  INV_X1    g013(.A(G197gat), .ZN(new_n215_));
  INV_X1    g014(.A(G204gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G197gat), .A2(G204gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n210_), .B1(KEYINPUT93), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n212_), .A2(new_n214_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G141gat), .ZN(new_n224_));
  INV_X1    g023(.A(G148gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n224_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT90), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT90), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(new_n224_), .A3(new_n225_), .A4(KEYINPUT90), .ZN(new_n230_));
  AND3_X1   g029(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT89), .B1(new_n235_), .B2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT1), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT88), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(G141gat), .B2(G148gat), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n246_), .A2(new_n248_), .B1(G141gat), .B2(G148gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n238_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n205_), .B(new_n223_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n219_), .A2(KEYINPUT93), .ZN(new_n254_));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n222_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n209_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n213_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n238_), .A2(new_n250_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n253_), .B1(new_n205_), .B2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G78gat), .B(G106gat), .Z(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n264_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n251_), .A2(new_n252_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n268_), .B(KEYINPUT28), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n271_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n275_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G8gat), .B(G36gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G183gat), .ZN(new_n286_));
  INV_X1    g085(.A(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT81), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT23), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT23), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT95), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT95), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G169gat), .A3(G176gat), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n298_), .A2(new_n299_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n299_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n306_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n292_), .A2(KEYINPUT23), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n290_), .A2(KEYINPUT81), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n289_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n295_), .A2(new_n290_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n286_), .A2(KEYINPUT25), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G183gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n287_), .A2(KEYINPUT26), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G190gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .A4(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n305_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n323_), .B2(new_n223_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n288_), .B(new_n314_), .C1(new_n325_), .C2(new_n295_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT83), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n313_), .A2(new_n328_), .A3(new_n288_), .A4(new_n314_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n300_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n308_), .A2(KEYINPUT22), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n308_), .A2(KEYINPUT22), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT82), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n308_), .A2(KEYINPUT22), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  AOI21_X1  g134(.A(G176gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n327_), .A2(new_n329_), .A3(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n294_), .A2(new_n296_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n318_), .A2(new_n320_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n315_), .A2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n315_), .A2(new_n317_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n340_), .B(new_n342_), .C1(new_n343_), .C2(new_n341_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n344_), .A3(new_n310_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n259_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT19), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n324_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT20), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n323_), .B2(new_n223_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n259_), .A3(new_n345_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n285_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n348_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n338_), .A2(new_n345_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n223_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n313_), .A2(new_n321_), .A3(new_n314_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n360_), .A2(new_n310_), .B1(new_n297_), .B2(new_n304_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n351_), .B1(new_n361_), .B2(new_n259_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n362_), .A3(new_n350_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n284_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(new_n364_), .A3(KEYINPUT96), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n357_), .A2(new_n363_), .A3(new_n366_), .A4(new_n284_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT105), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT105), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n365_), .A2(new_n371_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n348_), .B1(new_n324_), .B2(new_n346_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n352_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n284_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n377_), .A2(KEYINPUT27), .A3(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT106), .B1(new_n373_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT106), .ZN(new_n381_));
  AOI211_X1 g180(.A(new_n381_), .B(new_n378_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n280_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G127gat), .B(G134gat), .Z(new_n384_));
  XOR2_X1   g183(.A(G113gat), .B(G120gat), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n260_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n238_), .A2(new_n250_), .A3(new_n390_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT4), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT97), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT98), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n390_), .B1(new_n238_), .B2(new_n250_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n394_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n395_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT102), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G85gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT100), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT100), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n392_), .A2(new_n413_), .A3(new_n393_), .A4(new_n397_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n405_), .A2(new_n406_), .A3(new_n410_), .A4(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n238_), .A2(new_n250_), .A3(new_n390_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n417_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n260_), .A2(new_n391_), .A3(new_n401_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n398_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT99), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n394_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n415_), .A2(new_n421_), .A3(new_n410_), .A4(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT102), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n415_), .A2(new_n422_), .A3(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n410_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n416_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT103), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n416_), .A2(new_n424_), .A3(KEYINPUT103), .A4(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n434_), .A2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(G15gat), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G227gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n202_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n434_), .A2(new_n435_), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n436_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n441_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT84), .B(G43gat), .Z(new_n447_));
  NOR3_X1   g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n437_), .A2(G15gat), .A3(new_n438_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n443_), .B1(new_n442_), .B2(new_n436_), .ZN(new_n451_));
  OAI22_X1  g250(.A1(new_n450_), .A2(new_n451_), .B1(new_n440_), .B2(new_n202_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n439_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n358_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n338_), .A2(KEYINPUT30), .A3(new_n345_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT86), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(KEYINPUT86), .A3(new_n458_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n455_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n447_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(new_n449_), .A3(new_n453_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n459_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT31), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n461_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n469_), .B2(new_n459_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT87), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n391_), .A3(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n467_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n390_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n433_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n374_), .A2(new_n375_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n284_), .A2(KEYINPUT32), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n482_), .A2(KEYINPUT101), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n357_), .A2(new_n363_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT101), .B1(new_n486_), .B2(new_n483_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n484_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n428_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n365_), .A2(new_n367_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n394_), .A2(new_n397_), .A3(new_n419_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n392_), .A2(new_n393_), .A3(new_n398_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n491_), .A2(new_n426_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n423_), .B2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n490_), .B(new_n495_), .C1(new_n494_), .C2(new_n423_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n279_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n430_), .A2(new_n279_), .A3(new_n431_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n378_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n480_), .A2(new_n477_), .ZN(new_n501_));
  OAI22_X1  g300(.A1(new_n383_), .A2(new_n481_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT77), .B(G15gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G22gat), .ZN(new_n504_));
  INV_X1    g303(.A(G1gat), .ZN(new_n505_));
  INV_X1    g304(.A(G8gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G1gat), .B(G8gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n510_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT78), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(G229gat), .A3(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n513_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n516_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G169gat), .B(G197gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(KEYINPUT79), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n516_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n523_), .A2(new_n526_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n502_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT107), .Z(new_n535_));
  XOR2_X1   g334(.A(G120gat), .B(G148gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT71), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT6), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT65), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(G85gat), .ZN(new_n547_));
  INV_X1    g346(.A(G92gat), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT9), .ZN(new_n549_));
  XOR2_X1   g348(.A(G85gat), .B(G92gat), .Z(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(KEYINPUT9), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT10), .B(G99gat), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n546_), .B(new_n551_), .C1(G106gat), .C2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT8), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT7), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n546_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n544_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n555_), .B1(new_n560_), .B2(new_n550_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n554_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT67), .Z(new_n563_));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT68), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT11), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n566_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n570_), .A3(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n563_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n562_), .B(KEYINPUT67), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT64), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT69), .Z(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n575_), .A2(KEYINPUT12), .A3(new_n562_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n573_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT70), .B1(new_n585_), .B2(new_n579_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n573_), .A2(new_n584_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n588_));
  INV_X1    g387(.A(new_n579_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(new_n583_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n542_), .B1(new_n581_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n580_), .B(KEYINPUT69), .ZN(new_n593_));
  INV_X1    g392(.A(new_n542_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n586_), .A4(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n595_), .A3(KEYINPUT13), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n572_), .B(new_n510_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n604_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n563_), .A2(new_n513_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT74), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n618_), .B(new_n619_), .C1(new_n562_), .C2(new_n518_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(KEYINPUT74), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT73), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT36), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n627_), .B(KEYINPUT36), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n623_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n634_));
  AND3_X1   g433(.A1(new_n631_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n632_), .B(KEYINPUT75), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n623_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n631_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n600_), .A2(new_n613_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n535_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n505_), .A3(new_n432_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n598_), .A2(new_n599_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n613_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n502_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n631_), .A2(new_n633_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n647_), .A2(new_n533_), .A3(new_n648_), .A4(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n433_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n644_), .A2(new_n645_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n653_), .A3(new_n654_), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n380_), .A2(new_n382_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n643_), .A2(new_n506_), .A3(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT108), .Z(new_n658_));
  INV_X1    g457(.A(new_n656_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n652_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n506_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n661_), .B2(new_n660_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n662_), .B(KEYINPUT39), .C1(new_n661_), .C2(new_n660_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n658_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n658_), .B2(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  NAND3_X1  g470(.A1(new_n643_), .A2(new_n443_), .A3(new_n501_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n480_), .A2(new_n477_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G15gat), .B1(new_n652_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT41), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n674_), .A3(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n652_), .B2(new_n280_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n280_), .A2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n642_), .B2(new_n681_), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n650_), .A2(new_n613_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n600_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n535_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n432_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n635_), .A2(new_n639_), .A3(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n649_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n502_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n373_), .A2(new_n379_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n430_), .A2(new_n279_), .A3(new_n431_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n675_), .B1(new_n695_), .B2(new_n497_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(KEYINPUT112), .C1(new_n383_), .C2(new_n481_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n640_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n690_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n598_), .A2(new_n533_), .A3(new_n599_), .A4(new_n613_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT111), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n688_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n698_), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT113), .B1(new_n698_), .B2(KEYINPUT43), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n707_), .A2(new_n708_), .B1(new_n649_), .B2(new_n689_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n704_), .B(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(KEYINPUT44), .A3(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n432_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n687_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n685_), .A2(G36gat), .A3(new_n659_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT45), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n656_), .A3(new_n712_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G36gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT46), .B(new_n717_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  NAND4_X1  g525(.A1(new_n706_), .A2(G43gat), .A3(new_n712_), .A4(new_n501_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT115), .ZN(new_n728_));
  INV_X1    g527(.A(G43gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n685_), .B2(new_n675_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(KEYINPUT115), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n728_), .A2(new_n734_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n686_), .B2(new_n279_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n279_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n713_), .B2(new_n738_), .ZN(G1331gat));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n649_), .A2(new_n533_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n640_), .A2(new_n613_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n600_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n743_), .B2(new_n433_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT116), .ZN(new_n745_));
  INV_X1    g544(.A(new_n533_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n651_), .A2(new_n600_), .A3(new_n746_), .A4(new_n648_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n740_), .A3(new_n433_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1332gat));
  OAI21_X1  g548(.A(G64gat), .B1(new_n747_), .B2(new_n659_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT48), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n659_), .A2(G64gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n743_), .B2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n747_), .B2(new_n675_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n675_), .A2(G71gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n743_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT117), .Z(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n747_), .B2(new_n280_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n280_), .A2(G78gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n743_), .B2(new_n762_), .ZN(G1335gat));
  NAND4_X1  g562(.A1(new_n741_), .A2(new_n600_), .A3(new_n613_), .A4(new_n650_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n547_), .B1(new_n764_), .B2(new_n433_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT119), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n647_), .A2(new_n533_), .A3(new_n648_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n709_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n433_), .A2(new_n547_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NOR3_X1   g570(.A1(new_n764_), .A2(G92gat), .A3(new_n659_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n656_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G92gat), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT120), .ZN(G1337gat));
  NAND2_X1  g574(.A1(new_n501_), .A2(new_n552_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI22_X1  g576(.A1(new_n764_), .A2(new_n776_), .B1(KEYINPUT121), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n769_), .A2(new_n501_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G99gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(KEYINPUT121), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n780_), .B(new_n781_), .Z(G1338gat));
  XNOR2_X1  g581(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n709_), .A2(new_n279_), .A3(new_n767_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n764_), .A2(G106gat), .A3(new_n280_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n783_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n789_), .B(new_n783_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n647_), .A2(new_n746_), .A3(new_n742_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT54), .Z(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n585_), .A2(new_n797_), .A3(new_n579_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n589_), .B1(new_n587_), .B2(new_n583_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n586_), .A2(new_n590_), .A3(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n540_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n541_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n515_), .A2(new_n520_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n520_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n526_), .B1(new_n519_), .B2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n527_), .A2(new_n530_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n593_), .A2(new_n541_), .A3(new_n586_), .A4(new_n590_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n796_), .B1(new_n806_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n812_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(KEYINPUT58), .C1(new_n803_), .C2(new_n805_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n815_), .A3(new_n640_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n533_), .B(new_n811_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n596_), .A2(new_n810_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n650_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(KEYINPUT57), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT123), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n816_), .B(new_n822_), .C1(KEYINPUT57), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n795_), .B1(new_n825_), .B2(new_n613_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n383_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n675_), .A2(new_n433_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT124), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n833_));
  INV_X1    g632(.A(new_n824_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n820_), .B2(KEYINPUT123), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n648_), .B1(new_n835_), .B2(new_n823_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n833_), .B(new_n830_), .C1(new_n836_), .C2(new_n795_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n613_), .B1(new_n820_), .B2(new_n834_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n794_), .B(KEYINPUT54), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n829_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n832_), .A2(new_n533_), .A3(new_n837_), .A4(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G113gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n829_), .ZN(new_n844_));
  INV_X1    g643(.A(G113gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n533_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1340gat));
  NAND4_X1  g646(.A1(new_n832_), .A2(new_n600_), .A3(new_n837_), .A4(new_n841_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G120gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n838_), .A2(new_n839_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  AOI21_X1  g650(.A(G120gat), .B1(new_n600_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n851_), .B2(G120gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n850_), .A2(new_n827_), .A3(new_n828_), .A4(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT125), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n849_), .A2(new_n855_), .ZN(G1341gat));
  NAND4_X1  g655(.A1(new_n832_), .A2(new_n648_), .A3(new_n837_), .A4(new_n841_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G127gat), .ZN(new_n858_));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n844_), .A2(new_n859_), .A3(new_n648_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1342gat));
  NAND4_X1  g660(.A1(new_n832_), .A2(new_n640_), .A3(new_n837_), .A4(new_n841_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G134gat), .ZN(new_n863_));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n844_), .A2(new_n864_), .A3(new_n650_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n840_), .A2(new_n501_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n656_), .A2(new_n280_), .A3(new_n433_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n224_), .A3(new_n533_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G141gat), .B1(new_n869_), .B2(new_n746_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1344gat));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n225_), .A3(new_n600_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G148gat), .B1(new_n869_), .B2(new_n647_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1345gat));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n869_), .A2(new_n613_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n613_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(new_n640_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G162gat), .B1(new_n869_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n650_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n869_), .B2(new_n884_), .ZN(G1347gat));
  NOR3_X1   g684(.A1(new_n659_), .A2(new_n279_), .A3(new_n481_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n533_), .B(new_n886_), .C1(new_n836_), .C2(new_n795_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G169gat), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n298_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n890_), .B(new_n891_), .C1(new_n892_), .C2(new_n887_), .ZN(G1348gat));
  NOR2_X1   g692(.A1(new_n659_), .A2(new_n481_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n600_), .A2(G176gat), .A3(new_n894_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n840_), .A2(new_n279_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n826_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n600_), .A3(new_n886_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n299_), .ZN(G1349gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n886_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n900_), .A2(new_n343_), .A3(new_n613_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n850_), .A2(new_n280_), .A3(new_n648_), .A4(new_n894_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n902_), .A2(new_n286_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1350gat));
  OAI211_X1 g703(.A(new_n640_), .B(new_n886_), .C1(new_n836_), .C2(new_n795_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n905_), .A2(new_n906_), .A3(G190gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n905_), .B2(G190gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n650_), .A2(new_n340_), .ZN(new_n909_));
  OAI22_X1  g708(.A1(new_n907_), .A2(new_n908_), .B1(new_n900_), .B2(new_n909_), .ZN(G1351gat));
  NOR2_X1   g709(.A1(new_n659_), .A2(new_n694_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n867_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912_), .B2(new_n533_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n867_), .A2(new_n911_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n914_), .A2(new_n215_), .A3(new_n746_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1352gat));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n216_), .A3(new_n600_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G204gat), .B1(new_n914_), .B2(new_n647_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1353gat));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n648_), .A3(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n914_), .B2(new_n613_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n912_), .A2(new_n925_), .A3(new_n650_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G218gat), .B1(new_n914_), .B2(new_n881_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1355gat));
endmodule


