//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n209_), .B(new_n210_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n202_), .B1(new_n205_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n202_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n208_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n216_), .A2(new_n212_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G22gat), .B(G50gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT28), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n222_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(G211gat), .B(G218gat), .Z(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT21), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n226_), .A3(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(KEYINPUT88), .A3(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n221_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(G228gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n234_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n244_), .B1(new_n247_), .B2(new_n239_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G78gat), .B(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n225_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(KEYINPUT89), .A3(new_n250_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n253_), .A3(new_n225_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT89), .B1(new_n249_), .B2(new_n250_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT90), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n253_), .A2(new_n225_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .A4(new_n255_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n254_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT91), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT91), .ZN(new_n270_));
  AOI21_X1  g069(.A(G176gat), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n274_), .B(new_n275_), .C1(G183gat), .C2(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n282_), .A2(G169gat), .A3(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT82), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n281_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT25), .B(G183gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n274_), .A2(new_n275_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT82), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n282_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT24), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(G169gat), .B2(G176gat), .ZN(new_n297_));
  OAI22_X1  g096(.A1(new_n271_), .A2(new_n280_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n267_), .B1(new_n298_), .B2(new_n234_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n284_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT22), .B1(new_n284_), .B2(KEYINPUT84), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n285_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n276_), .B(new_n279_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n277_), .B(KEYINPUT83), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(new_n296_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n293_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n236_), .A2(new_n307_), .A3(new_n237_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n266_), .B1(new_n299_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n238_), .A2(new_n306_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n269_), .A2(new_n270_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n285_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n280_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n293_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n297_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n313_), .A2(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n267_), .B1(new_n317_), .B2(new_n247_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n318_), .A3(new_n266_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G64gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G92gat), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n310_), .B(new_n319_), .C1(new_n320_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n266_), .B1(new_n311_), .B2(new_n318_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n299_), .A2(new_n308_), .A3(new_n266_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT32), .B(new_n326_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G57gat), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n214_), .A2(new_n219_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G127gat), .B(G134gat), .Z(new_n337_));
  XOR2_X1   g136(.A(G113gat), .B(G120gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n214_), .A3(new_n219_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT4), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n336_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n335_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n335_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n334_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n346_), .A2(new_n334_), .A3(new_n348_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n325_), .B(new_n329_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n310_), .A2(new_n326_), .A3(new_n319_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n334_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n341_), .A2(new_n342_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n347_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT33), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n347_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n354_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n343_), .A2(new_n345_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n347_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  INV_X1    g162(.A(new_n348_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n362_), .A2(KEYINPUT93), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n307_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n234_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n265_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n324_), .B1(new_n368_), .B2(new_n309_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n353_), .A2(new_n360_), .A3(new_n365_), .A4(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n349_), .B2(KEYINPUT93), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n352_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n263_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n306_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT30), .B(new_n303_), .C1(new_n293_), .C2(new_n305_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n375_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n379_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n279_), .A2(KEYINPUT24), .A3(new_n294_), .A4(new_n295_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n291_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n287_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT30), .B1(new_n387_), .B2(new_n303_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n378_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n384_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n374_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n382_), .A2(new_n383_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n383_), .B1(new_n382_), .B2(new_n392_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT31), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n382_), .A2(new_n392_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n383_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n394_), .A3(new_n393_), .A4(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n340_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n402_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n339_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n373_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n258_), .A2(new_n262_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n254_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n397_), .A2(new_n340_), .A3(new_n402_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n340_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n263_), .A3(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n353_), .A2(new_n369_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n353_), .A3(KEYINPUT27), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n350_), .A2(new_n351_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n406_), .B1(new_n414_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G127gat), .B(G155gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G183gat), .B(G211gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n428_), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT17), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n428_), .B(new_n429_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n432_), .A2(new_n435_), .A3(KEYINPUT79), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT79), .B1(new_n435_), .B2(new_n432_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(KEYINPUT11), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n443_));
  XOR2_X1   g242(.A(G71gat), .B(G78gat), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n439_), .A3(KEYINPUT11), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(KEYINPUT11), .B2(new_n440_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n441_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G8gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453_));
  INV_X1    g252(.A(G8gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT75), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n456_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(G8gat), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT14), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G15gat), .B(G22gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n453_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  AOI211_X1 g267(.A(KEYINPUT76), .B(new_n466_), .C1(new_n459_), .C2(new_n464_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n452_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n457_), .A2(KEYINPUT75), .A3(new_n458_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n463_), .B1(new_n462_), .B2(KEYINPUT14), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n467_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT76), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n453_), .A3(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n451_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G231gat), .ZN(new_n477_));
  INV_X1    g276(.A(G233gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n470_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n450_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n470_), .A2(new_n476_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n479_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n450_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n470_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n438_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n432_), .B(KEYINPUT78), .Z(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n425_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n438_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n483_), .A2(new_n488_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT80), .B(new_n493_), .C1(new_n494_), .C2(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT34), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT35), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT70), .ZN(new_n500_));
  XOR2_X1   g299(.A(G29gat), .B(G36gat), .Z(new_n501_));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n506_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(KEYINPUT64), .A3(new_n522_), .ZN(new_n526_));
  AOI21_X1  g325(.A(G106gat), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n513_), .A2(new_n529_), .A3(new_n514_), .ZN(new_n530_));
  OR3_X1    g329(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n510_), .A2(new_n511_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n508_), .A3(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  AND2_X1   g339(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n541_));
  NOR2_X1   g340(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(new_n543_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n515_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n536_), .B1(new_n546_), .B2(new_n529_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n528_), .B1(new_n547_), .B2(KEYINPUT68), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n529_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n549_), .A2(KEYINPUT68), .A3(new_n535_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n505_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n525_), .A2(new_n526_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n519_), .B1(new_n553_), .B2(G106gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n549_), .B2(new_n535_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n503_), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n555_), .A2(new_n556_), .B1(KEYINPUT35), .B2(new_n498_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n500_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n503_), .B(KEYINPUT15), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n549_), .A2(new_n535_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n554_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n500_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT36), .Z(new_n570_));
  NAND3_X1  g369(.A1(new_n558_), .A2(new_n566_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT72), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n558_), .A2(new_n573_), .A3(new_n566_), .A4(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n558_), .A2(new_n566_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(KEYINPUT36), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT71), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n579_), .A2(new_n580_), .A3(KEYINPUT37), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n579_), .B2(KEYINPUT37), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n571_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT37), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n581_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n424_), .A2(new_n496_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n450_), .A2(KEYINPUT12), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n563_), .B2(new_n550_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n555_), .A2(new_n450_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n561_), .A2(new_n528_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(new_n486_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n486_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n590_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  INV_X1    g400(.A(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT5), .B(G176gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n600_), .A2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n587_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n600_), .A2(new_n605_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT13), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n468_), .A2(new_n469_), .A3(new_n452_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n451_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n503_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n470_), .A2(new_n476_), .A3(new_n556_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n484_), .B2(new_n503_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n470_), .A2(new_n476_), .A3(new_n560_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n617_), .A2(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(new_n284_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(G197gat), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n470_), .A2(new_n476_), .A3(new_n556_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n556_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n619_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n615_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n625_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT81), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT81), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n629_), .A2(new_n630_), .A3(new_n633_), .A4(new_n625_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n626_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n612_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n586_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(KEYINPUT94), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n421_), .B(KEYINPUT95), .Z(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n461_), .A3(new_n460_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(new_n641_), .A3(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n637_), .B(new_n639_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n489_), .A2(new_n491_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n612_), .A2(new_n635_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n414_), .A2(new_n423_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n406_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n658_), .A3(new_n583_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n421_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n648_), .A2(new_n650_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n648_), .A2(new_n650_), .A3(KEYINPUT98), .A4(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n454_), .A3(new_n420_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668_));
  INV_X1    g467(.A(new_n420_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n659_), .B2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(G8gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n659_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT99), .A3(new_n420_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n667_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  AND4_X1   g473(.A1(new_n667_), .A2(new_n673_), .A3(G8gat), .A4(new_n670_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n666_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT40), .Z(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n666_), .B(new_n678_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1325gat));
  NOR2_X1   g481(.A1(new_n410_), .A2(new_n411_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G15gat), .B1(new_n659_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n637_), .A2(G15gat), .A3(new_n684_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(G1326gat));
  INV_X1    g489(.A(G22gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n409_), .B(KEYINPUT103), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n672_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT42), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n638_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n496_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n583_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n658_), .A2(KEYINPUT105), .A3(new_n636_), .A4(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n423_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n636_), .B(new_n698_), .C1(new_n701_), .C2(new_n406_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n422_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n579_), .A2(KEYINPUT37), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT73), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n579_), .A2(new_n580_), .A3(KEYINPUT37), .ZN(new_n711_));
  INV_X1    g510(.A(new_n584_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n424_), .B2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT43), .B(new_n585_), .C1(new_n701_), .C2(new_n406_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(new_n636_), .A3(new_n496_), .A4(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT104), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n642_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n707_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n721_), .B2(new_n420_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n669_), .A2(G36gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n699_), .A2(new_n704_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT106), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n699_), .A2(new_n704_), .A3(new_n730_), .A4(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(KEYINPUT45), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n724_), .B1(new_n726_), .B2(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n716_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n716_), .B2(KEYINPUT104), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n420_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT46), .A3(new_n735_), .A4(new_n734_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1329gat));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n683_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G43gat), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n705_), .A2(G43gat), .A3(new_n684_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT47), .B(new_n747_), .C1(new_n745_), .C2(G43gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n706_), .B2(new_n692_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n409_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n721_), .B2(new_n753_), .ZN(G1331gat));
  INV_X1    g553(.A(new_n583_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n424_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n612_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n632_), .A2(new_n634_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n622_), .A2(new_n625_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n492_), .A2(new_n495_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n421_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n759_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n757_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n586_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n643_), .A2(G57gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g568(.A(G64gat), .B1(new_n762_), .B2(new_n669_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT48), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n669_), .A2(G64gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n766_), .B2(new_n772_), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n762_), .B2(new_n684_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n684_), .A2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n766_), .B2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  INV_X1    g577(.A(new_n762_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n692_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT50), .Z(new_n781_));
  NAND2_X1  g580(.A1(new_n692_), .A2(new_n778_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n766_), .B2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n424_), .A2(new_n697_), .A3(new_n583_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n765_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n642_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n714_), .A2(new_n496_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n715_), .A3(new_n765_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n422_), .A2(G85gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT108), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n787_), .B1(new_n790_), .B2(new_n792_), .ZN(G1336gat));
  OAI21_X1  g592(.A(G92gat), .B1(new_n789_), .B2(new_n669_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n785_), .A2(G92gat), .A3(new_n669_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT109), .Z(G1337gat));
  OR3_X1    g596(.A1(new_n785_), .A2(new_n553_), .A3(new_n684_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n788_), .A2(new_n683_), .A3(new_n715_), .A4(new_n765_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(G99gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G99gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT51), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n798_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1338gat));
  OR3_X1    g606(.A1(new_n785_), .A2(G106gat), .A3(new_n263_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n788_), .A2(new_n409_), .A3(new_n715_), .A4(new_n765_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G106gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G106gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n814_), .B(new_n808_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n589_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n593_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n822_));
  NAND2_X1  g621(.A1(new_n596_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .A4(KEYINPUT55), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n605_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n608_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n610_), .A2(new_n606_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n615_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n625_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n632_), .A2(new_n634_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n830_), .A2(new_n831_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n836_), .A2(new_n755_), .B1(new_n837_), .B2(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n764_), .A2(new_n610_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n605_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n583_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n835_), .B(new_n610_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n835_), .A2(new_n610_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n830_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n850_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n585_), .A2(new_n851_), .A3(new_n853_), .A4(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n651_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n760_), .A2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n635_), .A2(KEYINPUT112), .A3(new_n492_), .A4(new_n495_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n757_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n860_), .B2(new_n585_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n859_), .A2(new_n757_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n713_), .A4(new_n858_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n819_), .B1(new_n856_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n864_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n851_), .A2(new_n853_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT58), .B1(new_n852_), .B2(new_n830_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n713_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n870_), .B1(new_n838_), .B2(new_n846_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT116), .B(new_n867_), .C1(new_n871_), .C2(new_n651_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n413_), .A2(new_n643_), .A3(new_n420_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G113gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n764_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n847_), .A2(new_n855_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n496_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n881_), .B2(new_n867_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n635_), .B(new_n882_), .C1(new_n874_), .C2(KEYINPUT59), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n877_), .B1(new_n883_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g683(.A(G120gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT60), .B1(new_n612_), .B2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(KEYINPUT60), .B2(new_n885_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n875_), .A2(KEYINPUT118), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT118), .B1(new_n875_), .B2(new_n887_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n757_), .B(new_n882_), .C1(new_n874_), .C2(KEYINPUT59), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n890_), .B2(new_n885_), .ZN(G1341gat));
  INV_X1    g690(.A(G127gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n875_), .A2(new_n892_), .A3(new_n697_), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n652_), .B(new_n882_), .C1(new_n874_), .C2(KEYINPUT59), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n892_), .ZN(G1342gat));
  INV_X1    g694(.A(G134gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n875_), .A2(new_n896_), .A3(new_n755_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n713_), .B(new_n882_), .C1(new_n874_), .C2(KEYINPUT59), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1343gat));
  AND2_X1   g698(.A1(new_n866_), .A2(new_n872_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n684_), .A2(new_n409_), .A3(new_n669_), .A4(new_n642_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n635_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n207_), .ZN(G1344gat));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n757_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n208_), .ZN(G1345gat));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n496_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT61), .B(G155gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n903_), .B2(new_n713_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n583_), .A2(G162gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n903_), .B2(new_n912_), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n881_), .A2(new_n867_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n643_), .A2(new_n683_), .A3(new_n420_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n692_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n764_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT119), .B(KEYINPUT62), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n919_), .A2(G169gat), .A3(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n918_), .A2(new_n764_), .A3(new_n312_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n919_), .B2(G169gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n915_), .A2(new_n409_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n900_), .A2(G176gat), .A3(new_n612_), .A4(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n914_), .A2(new_n612_), .A3(new_n916_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n926_), .A2(new_n927_), .B1(new_n285_), .B2(new_n929_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n900_), .A2(new_n697_), .A3(new_n925_), .ZN(new_n932_));
  INV_X1    g731(.A(G183gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n652_), .A2(new_n288_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n932_), .A2(new_n933_), .B1(new_n918_), .B2(new_n934_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n917_), .B2(new_n713_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n755_), .A2(new_n289_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT121), .Z(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n917_), .B2(new_n938_), .ZN(G1351gat));
  OR2_X1    g738(.A1(new_n412_), .A2(new_n422_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n420_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n941_), .B2(new_n940_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n866_), .A2(new_n872_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n764_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g745(.A1(new_n866_), .A2(new_n872_), .A3(new_n612_), .A4(new_n943_), .ZN(new_n947_));
  OR3_X1    g746(.A1(new_n947_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n947_), .B2(G204gat), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n944_), .A2(new_n951_), .A3(new_n612_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n602_), .B1(new_n947_), .B2(KEYINPUT123), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n952_), .A2(new_n953_), .A3(KEYINPUT124), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT124), .B1(new_n952_), .B2(new_n953_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n950_), .B1(new_n954_), .B2(new_n955_), .ZN(G1353gat));
  AOI21_X1  g755(.A(new_n652_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n866_), .A2(new_n872_), .A3(new_n943_), .A4(new_n957_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n958_), .A2(KEYINPUT126), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(KEYINPUT126), .ZN(new_n960_));
  OR2_X1    g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  OR3_X1    g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n959_), .B2(new_n960_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1354gat));
  NAND4_X1  g763(.A1(new_n866_), .A2(new_n872_), .A3(new_n585_), .A4(new_n943_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(G218gat), .ZN(new_n966_));
  INV_X1    g765(.A(new_n944_), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n583_), .A2(G218gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(KEYINPUT127), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971_));
  OAI211_X1 g770(.A(new_n971_), .B(new_n966_), .C1(new_n967_), .C2(new_n968_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n972_), .ZN(G1355gat));
endmodule


