//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT77), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT68), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n208_), .A2(KEYINPUT68), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(KEYINPUT68), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n210_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT76), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT74), .B(G8gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G1gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G1gat), .B(G8gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n207_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(new_n218_), .A3(KEYINPUT77), .A4(new_n220_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n216_), .B(new_n233_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n230_), .A2(new_n232_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n231_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n239_));
  AOI211_X1 g038(.A(new_n236_), .B(new_n239_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n206_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n237_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n205_), .C1(new_n237_), .C2(new_n235_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G141gat), .ZN(new_n246_));
  INV_X1    g045(.A(G148gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT85), .B1(new_n248_), .B2(KEYINPUT3), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT86), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  AND2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n262_), .A2(KEYINPUT1), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT83), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n262_), .A2(new_n275_), .A3(KEYINPUT1), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n246_), .A2(new_n247_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n250_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(KEYINPUT84), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT84), .B1(new_n277_), .B2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n270_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n282_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n268_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n261_), .B1(KEYINPUT1), .B2(new_n262_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n262_), .A2(new_n275_), .A3(KEYINPUT1), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n275_), .B1(new_n262_), .B2(KEYINPUT1), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n279_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n285_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n277_), .A2(KEYINPUT84), .A3(new_n279_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT28), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n283_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G22gat), .B(G50gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n283_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT88), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n291_), .A2(new_n292_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n294_), .B1(new_n306_), .B2(new_n270_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT21), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  INV_X1    g112(.A(new_n309_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n305_), .B1(new_n307_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n282_), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n318_), .A2(new_n305_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT87), .B1(new_n282_), .B2(KEYINPUT29), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n328_), .A2(KEYINPUT89), .A3(new_n322_), .A4(new_n323_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n320_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT90), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n302_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n329_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n319_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n337_), .A3(KEYINPUT91), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT91), .ZN(new_n339_));
  INV_X1    g138(.A(new_n323_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n307_), .B2(KEYINPUT87), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT89), .B1(new_n341_), .B2(new_n328_), .ZN(new_n342_));
  AND4_X1   g141(.A1(KEYINPUT89), .A2(new_n328_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n319_), .B(new_n332_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n301_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n298_), .B1(new_n283_), .B2(new_n296_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n332_), .B1(new_n334_), .B2(new_n319_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n334_), .A2(new_n319_), .A3(new_n331_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n302_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n330_), .A2(new_n331_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n338_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  NOR2_X1   g157(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n360_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(KEYINPUT81), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(new_n363_), .A3(G183gat), .A4(G190gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n361_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT80), .B1(new_n361_), .B2(KEYINPUT23), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n369_), .B(new_n371_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT25), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G183gat), .ZN(new_n379_));
  INV_X1    g178(.A(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT26), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT26), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G190gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n377_), .A2(new_n379_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n386_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n384_), .A2(new_n389_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n368_), .B1(new_n375_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n312_), .A2(new_n317_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT20), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n386_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT92), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n384_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n365_), .A2(new_n393_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n367_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n374_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n360_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n318_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n358_), .B1(new_n397_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n409_), .A3(new_n318_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n395_), .A2(new_n396_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n358_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT20), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(KEYINPUT93), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT18), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT25), .B(G183gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G190gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n392_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n374_), .A2(new_n423_), .A3(new_n391_), .A4(new_n389_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n318_), .A2(new_n424_), .A3(new_n368_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n421_), .A2(new_n422_), .B1(new_n398_), .B2(new_n386_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n404_), .B1(new_n426_), .B2(new_n402_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n427_), .A2(new_n401_), .B1(new_n408_), .B2(new_n360_), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT20), .B(new_n425_), .C1(new_n428_), .C2(new_n318_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n358_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n416_), .A2(new_n420_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n420_), .B1(new_n416_), .B2(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n356_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n416_), .A2(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n420_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT96), .B1(new_n429_), .B2(new_n358_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n397_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n406_), .A2(new_n409_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n396_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .A4(new_n414_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT20), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n358_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n420_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n447_), .A3(KEYINPUT27), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n434_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT98), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n434_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G127gat), .B(G134gat), .Z(new_n454_));
  XOR2_X1   g253(.A(G113gat), .B(G120gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n282_), .A2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n270_), .B(new_n456_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT4), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT94), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n458_), .A2(new_n462_), .A3(KEYINPUT4), .A4(new_n459_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n456_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G29gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(G85gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT0), .B(G57gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n458_), .A2(new_n459_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(new_n468_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n469_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n464_), .B1(new_n460_), .B2(KEYINPUT94), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n467_), .B1(new_n479_), .B2(new_n463_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n480_), .B2(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G71gat), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n395_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(new_n456_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT82), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT30), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT31), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n488_), .B(new_n492_), .Z(new_n493_));
  NOR2_X1   g292(.A1(new_n482_), .A2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n355_), .A2(new_n453_), .A3(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n478_), .A2(new_n434_), .A3(new_n448_), .A4(new_n481_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n338_), .C1(new_n350_), .C2(new_n354_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n348_), .A2(new_n339_), .A3(new_n349_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n352_), .A2(new_n353_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT91), .B1(new_n333_), .B2(new_n337_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n446_), .A2(KEYINPUT32), .A3(new_n436_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n435_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT95), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n435_), .A2(new_n506_), .A3(new_n503_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n502_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n482_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n461_), .A2(new_n467_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n473_), .B1(new_n475_), .B2(new_n468_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n416_), .A2(new_n420_), .A3(new_n431_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n512_), .A2(new_n437_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT33), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n476_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n474_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT33), .B(new_n473_), .C1(new_n480_), .C2(new_n476_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n493_), .B(new_n497_), .C1(new_n501_), .C2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n495_), .B1(new_n521_), .B2(KEYINPUT97), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n355_), .A2(new_n509_), .A3(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n493_), .A4(new_n497_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n245_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528_));
  XOR2_X1   g327(.A(G85gat), .B(G92gat), .Z(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT6), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT8), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(KEYINPUT64), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n536_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT64), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n532_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n529_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n539_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n543_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT10), .B(G99gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(G106gat), .ZN(new_n551_));
  INV_X1    g350(.A(G85gat), .ZN(new_n552_));
  INV_X1    g351(.A(G92gat), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT9), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n549_), .A2(new_n551_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n234_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n217_), .A2(new_n548_), .A3(new_n556_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n559_), .A3(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n558_), .A2(new_n569_), .A3(new_n559_), .A4(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT69), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT36), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n528_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT71), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n575_), .B(KEYINPUT36), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT72), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n571_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n527_), .B1(new_n584_), .B2(KEYINPUT37), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  INV_X1    g385(.A(new_n581_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n571_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n580_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT73), .B(new_n586_), .C1(new_n580_), .C2(new_n583_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT11), .ZN(new_n595_));
  XOR2_X1   g394(.A(G71gat), .B(G78gat), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n594_), .A2(KEYINPUT11), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT65), .B(KEYINPUT12), .Z(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n600_), .ZN(new_n604_));
  OR2_X1    g403(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n605_));
  INV_X1    g404(.A(new_n532_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n543_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n541_), .A2(new_n542_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n609_), .A2(new_n546_), .B1(KEYINPUT8), .B2(new_n538_), .ZN(new_n610_));
  AND4_X1   g409(.A1(new_n549_), .A2(new_n551_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n604_), .B(new_n605_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n548_), .A2(new_n556_), .A3(new_n600_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT66), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n603_), .B(new_n612_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT5), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n613_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n601_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n618_), .B(new_n623_), .C1(new_n615_), .C2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n617_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n625_), .A2(new_n615_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n622_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT13), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT13), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XOR2_X1   g439(.A(G183gat), .B(G211gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n600_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(new_n229_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT17), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n646_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(KEYINPUT75), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT75), .B(new_n645_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n593_), .A2(new_n638_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n526_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n224_), .A3(new_n482_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n638_), .A2(new_n245_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n654_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT99), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n580_), .A2(new_n588_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT100), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n482_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n658_), .A2(new_n659_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n660_), .A2(new_n671_), .A3(new_n672_), .ZN(G1324gat));
  INV_X1    g472(.A(new_n453_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n664_), .A2(new_n668_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G8gat), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n223_), .A3(new_n674_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1325gat));
  OAI21_X1  g482(.A(G15gat), .B1(new_n669_), .B2(new_n493_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT103), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n686_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n656_), .A2(G15gat), .A3(new_n493_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n669_), .B2(new_n355_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT42), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n355_), .A2(G22gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n656_), .B2(new_n693_), .ZN(G1327gat));
  NOR3_X1   g493(.A1(new_n638_), .A2(new_n245_), .A3(new_n662_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n591_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT43), .B(new_n696_), .C1(new_n522_), .C2(new_n525_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n501_), .A2(new_n520_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n497_), .A2(new_n493_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT97), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n495_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n525_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n698_), .B1(new_n703_), .B2(new_n593_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n695_), .B1(new_n697_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n695_), .C1(new_n697_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n670_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n580_), .A2(new_n588_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n654_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT104), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n638_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(new_n526_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n670_), .A2(G29gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT105), .Z(new_n718_));
  OAI21_X1  g517(.A(new_n710_), .B1(new_n716_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT106), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT106), .ZN(new_n722_));
  OAI21_X1  g521(.A(G36gat), .B1(new_n709_), .B2(new_n453_), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n715_), .A2(new_n724_), .A3(new_n674_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n721_), .B(new_n722_), .C1(new_n723_), .C2(new_n726_), .ZN(new_n727_));
  AND4_X1   g526(.A1(KEYINPUT106), .A2(new_n723_), .A3(new_n720_), .A4(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(new_n493_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(G43gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n707_), .A2(new_n708_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n707_), .A2(KEYINPUT107), .A3(new_n708_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G43gat), .B1(new_n715_), .B2(new_n730_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT108), .Z(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT47), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n709_), .A2(new_n744_), .A3(new_n355_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G50gat), .B1(new_n715_), .B2(new_n501_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n241_), .A2(new_n244_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n749_), .A2(new_n638_), .A3(new_n662_), .A4(new_n696_), .ZN(new_n750_));
  AOI211_X1 g549(.A(G57gat), .B(new_n670_), .C1(new_n750_), .C2(KEYINPUT109), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n750_), .A2(KEYINPUT109), .ZN(new_n752_));
  INV_X1    g551(.A(new_n638_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n245_), .A2(new_n662_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n668_), .A2(new_n482_), .A3(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n751_), .A2(new_n752_), .B1(G57gat), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT110), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n668_), .A2(new_n755_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G64gat), .B1(new_n759_), .B2(new_n453_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT48), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n453_), .A2(G64gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n750_), .B2(new_n762_), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n759_), .B2(new_n493_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT49), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n493_), .A2(G71gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n750_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT111), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n759_), .B2(new_n355_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n355_), .A2(G78gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n750_), .B2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n713_), .A2(new_n753_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n749_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n552_), .A3(new_n482_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n697_), .A2(new_n704_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n753_), .A2(new_n748_), .A3(new_n662_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n482_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n781_), .B2(new_n552_), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n775_), .A2(new_n553_), .A3(new_n674_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n674_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n553_), .ZN(G1337gat));
  OR3_X1    g585(.A1(new_n774_), .A2(new_n493_), .A3(new_n550_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n779_), .A2(new_n730_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n789_), .B2(new_n485_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT51), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n787_), .C1(new_n789_), .C2(new_n485_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1338gat));
  INV_X1    g593(.A(G106gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n775_), .A2(new_n795_), .A3(new_n501_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n501_), .A3(new_n778_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT113), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(KEYINPUT113), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n797_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n796_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n796_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  AOI21_X1  g606(.A(new_n206_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n241_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n626_), .B1(new_n811_), .B2(KEYINPUT58), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(KEYINPUT58), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n615_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n627_), .B2(new_n624_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n630_), .B2(KEYINPUT55), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n618_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n622_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n603_), .A2(new_n613_), .A3(new_n612_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n618_), .A2(new_n819_), .B1(new_n824_), .B2(new_n816_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n630_), .A2(KEYINPUT55), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n623_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT56), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n813_), .B(new_n815_), .C1(new_n823_), .C2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n813_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n814_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n593_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n748_), .A2(new_n626_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(KEYINPUT115), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n622_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n822_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n823_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n821_), .B2(KEYINPUT115), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n835_), .B1(new_n841_), .B2(new_n837_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n833_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n810_), .A2(new_n634_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n711_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n832_), .B1(new_n846_), .B2(KEYINPUT57), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n822_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n837_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n839_), .A3(new_n838_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n844_), .B1(new_n851_), .B2(new_n833_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n711_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n654_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n748_), .A2(new_n654_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n753_), .A2(KEYINPUT114), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n754_), .B2(new_n638_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n696_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n696_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n855_), .A2(new_n865_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n674_), .A2(new_n501_), .A3(new_n670_), .A4(new_n493_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n748_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n245_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n871_), .B1(new_n875_), .B2(new_n870_), .ZN(G1340gat));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n753_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n869_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n753_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n877_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n869_), .B2(new_n662_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n872_), .A2(new_n874_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n662_), .A2(G127gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT118), .Z(new_n885_));
  AOI21_X1  g684(.A(new_n882_), .B1(new_n883_), .B2(new_n885_), .ZN(G1342gat));
  AOI21_X1  g685(.A(G134gat), .B1(new_n869_), .B2(new_n667_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT119), .B(G134gat), .Z(new_n888_));
  NOR2_X1   g687(.A1(new_n696_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n883_), .B2(new_n889_), .ZN(G1343gat));
  XNOR2_X1  g689(.A(KEYINPUT121), .B(G141gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n355_), .B1(new_n855_), .B2(new_n865_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n674_), .A2(new_n670_), .A3(new_n730_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT120), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n896_), .A3(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n891_), .B1(new_n898_), .B2(new_n748_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n846_), .A2(KEYINPUT57), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n853_), .B1(new_n852_), .B2(new_n711_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n832_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n864_), .B1(new_n903_), .B2(new_n654_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n893_), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n904_), .A2(KEYINPUT120), .A3(new_n355_), .A4(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n748_), .B(new_n891_), .C1(new_n900_), .C2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n899_), .A2(new_n908_), .ZN(G1344gat));
  OAI21_X1  g708(.A(new_n638_), .B1(new_n900_), .B2(new_n906_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g710(.A(new_n662_), .B1(new_n900_), .B2(new_n906_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1346gat));
  INV_X1    g713(.A(G162gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n898_), .A2(new_n915_), .A3(new_n667_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n696_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(G1347gat));
  NAND2_X1  g717(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G169gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n674_), .A2(new_n494_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT122), .Z(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n355_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n904_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n920_), .B1(new_n924_), .B2(new_n748_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n926_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n866_), .A2(new_n929_), .A3(new_n355_), .A4(new_n922_), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT124), .B1(new_n904_), .B2(new_n923_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n748_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n927_), .A2(new_n928_), .B1(new_n932_), .B2(new_n935_), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n638_), .A2(new_n937_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n904_), .A2(new_n753_), .A3(new_n923_), .ZN(new_n939_));
  OAI22_X1  g738(.A1(new_n932_), .A2(new_n938_), .B1(new_n937_), .B2(new_n939_), .ZN(G1349gat));
  OR2_X1    g739(.A1(new_n654_), .A2(new_n421_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n942_));
  AOI21_X1  g741(.A(G183gat), .B1(new_n924_), .B2(new_n662_), .ZN(new_n943_));
  OR3_X1    g742(.A1(new_n942_), .A2(new_n943_), .A3(KEYINPUT125), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n943_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n932_), .B2(new_n696_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n667_), .A2(new_n422_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n932_), .B2(new_n948_), .ZN(G1351gat));
  NOR3_X1   g748(.A1(new_n453_), .A2(new_n482_), .A3(new_n730_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n892_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n748_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n638_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g754(.A(KEYINPUT63), .B(G211gat), .Z(new_n956_));
  AND3_X1   g755(.A1(new_n951_), .A2(new_n662_), .A3(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n951_), .A2(new_n662_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n958_), .B2(new_n959_), .ZN(G1354gat));
  XOR2_X1   g759(.A(KEYINPUT126), .B(G218gat), .Z(new_n961_));
  NAND4_X1  g760(.A1(new_n892_), .A2(new_n593_), .A3(new_n950_), .A4(new_n961_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n892_), .A2(new_n667_), .A3(new_n950_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n963_), .B2(new_n961_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(KEYINPUT127), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n966_), .B(new_n962_), .C1(new_n963_), .C2(new_n961_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(G1355gat));
endmodule


