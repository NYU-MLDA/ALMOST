//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  OR3_X1    g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT1), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n202_), .B2(new_n203_), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n204_), .B(new_n205_), .C1(G155gat), .C2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT85), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT84), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT3), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(new_n209_), .B2(KEYINPUT2), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n216_), .A3(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n211_), .B1(KEYINPUT84), .B2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223_));
  XOR2_X1   g022(.A(G155gat), .B(G162gat), .Z(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n213_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n228_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n234_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n213_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n213_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n222_), .A2(new_n224_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT86), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n245_), .B2(new_n225_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n236_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n240_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT4), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT4), .B1(new_n228_), .B2(new_n236_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n238_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n242_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n254_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G64gat), .B(G92gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G8gat), .B(G36gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266_));
  XOR2_X1   g065(.A(G197gat), .B(G204gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT87), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n267_), .A2(KEYINPUT21), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n268_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n271_), .A2(new_n272_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n268_), .B(new_n273_), .C1(new_n276_), .C2(new_n269_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  OR2_X1    g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT22), .B(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(G176gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT24), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT24), .A3(new_n283_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294_));
  OR3_X1    g093(.A1(new_n294_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n294_), .B2(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(G190gat), .ZN(new_n297_));
  AND4_X1   g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n288_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n278_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT90), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n293_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n280_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n288_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n275_), .A2(new_n277_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(KEYINPUT90), .A3(new_n306_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT20), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n305_), .A2(new_n306_), .A3(KEYINPUT89), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  INV_X1    g115(.A(new_n299_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n306_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT89), .B1(new_n305_), .B2(new_n306_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(new_n313_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n266_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT95), .B1(new_n314_), .B2(new_n321_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n300_), .A2(new_n307_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n312_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(new_n265_), .C1(new_n320_), .C2(new_n312_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n265_), .A2(new_n322_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n259_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n254_), .A2(KEYINPUT93), .A3(KEYINPUT33), .A4(new_n258_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n250_), .B1(KEYINPUT4), .B2(new_n248_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n241_), .B(new_n258_), .C1(new_n332_), .C2(new_n238_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n331_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n252_), .A2(new_n238_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n258_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n337_), .B(new_n338_), .C1(new_n238_), .C2(new_n248_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n309_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n312_), .B1(new_n342_), .B2(KEYINPUT20), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n320_), .A2(new_n313_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n264_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n264_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n314_), .A2(new_n321_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n347_), .A3(KEYINPUT92), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(new_n264_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n333_), .A2(KEYINPUT94), .A3(new_n334_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT94), .B1(new_n333_), .B2(new_n334_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n329_), .B1(new_n340_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n278_), .B1(new_n246_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G228gat), .A3(G233gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n278_), .C1(new_n246_), .C2(new_n357_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G78gat), .B(G106gat), .Z(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G22gat), .B(G50gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n246_), .B2(new_n357_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n246_), .A2(new_n366_), .A3(new_n357_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n365_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n371_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT88), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n359_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n373_), .B2(new_n370_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n364_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT88), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n372_), .B1(new_n371_), .B2(new_n367_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n368_), .A2(new_n369_), .A3(new_n365_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n364_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n379_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n236_), .B(KEYINPUT31), .Z(new_n387_));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT30), .B(G15gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n299_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G43gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n395_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n387_), .A2(new_n388_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n400_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n356_), .A2(new_n386_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n348_), .A2(new_n405_), .A3(new_n350_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n326_), .B1(new_n320_), .B2(new_n312_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n346_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n345_), .A2(KEYINPUT27), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(new_n259_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n364_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n383_), .A2(new_n377_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n375_), .B1(new_n382_), .B2(new_n381_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n399_), .A2(new_n402_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n384_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n415_), .B2(new_n384_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n404_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G57gat), .A2(G64gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G57gat), .A2(G64gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT11), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT11), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(G78gat), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n432_));
  INV_X1    g231(.A(G78gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n428_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n424_), .A2(new_n427_), .A3(new_n431_), .A4(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n426_), .B1(new_n425_), .B2(new_n421_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n429_), .A2(new_n430_), .A3(G78gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n433_), .B1(new_n432_), .B2(new_n428_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G231gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT75), .B(G15gat), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G22gat), .ZN(new_n444_));
  INV_X1    g243(.A(G1gat), .ZN(new_n445_));
  INV_X1    g244(.A(G8gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT14), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT75), .B(G15gat), .ZN(new_n448_));
  INV_X1    g247(.A(G22gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G8gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT76), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n451_), .B(new_n453_), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n442_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n456_));
  XNOR2_X1  g255(.A(G127gat), .B(G155gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G183gat), .B(G211gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT17), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n460_), .A2(KEYINPUT17), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n455_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(KEYINPUT78), .Z(new_n466_));
  XNOR2_X1  g265(.A(G134gat), .B(G162gat), .ZN(new_n467_));
  INV_X1    g266(.A(G218gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT72), .B(G190gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT36), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G92gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G85gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G92gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT8), .B1(new_n491_), .B2(KEYINPUT65), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n487_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT64), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(G92gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(G85gat), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n478_), .A2(KEYINPUT10), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n478_), .A2(KEYINPUT10), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n479_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n489_), .A2(G92gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n487_), .A2(G85gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT9), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n483_), .A2(new_n484_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n498_), .A2(new_n501_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n486_), .B(new_n491_), .C1(KEYINPUT65), .C2(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n494_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n476_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(KEYINPUT34), .Z(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n494_), .A2(new_n475_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n509_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n511_), .A2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n509_), .A2(new_n518_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n472_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n520_), .A2(KEYINPUT73), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n471_), .A2(KEYINPUT36), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n520_), .B2(KEYINPUT73), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT37), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n472_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(KEYINPUT74), .A3(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n523_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n466_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n420_), .A2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n435_), .A2(new_n439_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n508_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n440_), .A2(new_n506_), .A3(new_n494_), .A4(new_n507_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT67), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT67), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n508_), .A2(new_n548_), .A3(new_n538_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT68), .B1(new_n550_), .B2(new_n542_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n552_), .B(new_n543_), .C1(new_n547_), .C2(new_n549_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n545_), .B(new_n546_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G176gat), .B(G204gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n554_), .A2(new_n559_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n560_), .B(new_n561_), .C1(new_n562_), .C2(KEYINPUT13), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n560_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n451_), .B(new_n453_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(new_n475_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n475_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n454_), .A2(new_n476_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n475_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n568_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT79), .ZN(new_n578_));
  XOR2_X1   g377(.A(G169gat), .B(G197gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n573_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT80), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n567_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n537_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n445_), .A3(new_n259_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT38), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n333_), .A2(new_n334_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n352_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(new_n351_), .A3(new_n339_), .A4(new_n336_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n416_), .B1(new_n598_), .B2(new_n329_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n403_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n415_), .A2(new_n416_), .A3(new_n384_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n599_), .A2(new_n386_), .B1(new_n602_), .B2(new_n411_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n531_), .A2(new_n523_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n465_), .A3(new_n589_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n259_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n593_), .A2(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n410_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G8gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT97), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n615_), .A3(G8gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(KEYINPUT39), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n612_), .B2(G8gat), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT97), .B(new_n446_), .C1(new_n611_), .C2(new_n410_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n591_), .A2(new_n446_), .A3(new_n410_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n617_), .A2(new_n621_), .A3(KEYINPUT40), .A4(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n607_), .B2(new_n403_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n403_), .A2(G15gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n590_), .B2(new_n631_), .ZN(G1326gat));
  OAI21_X1  g431(.A(G22gat), .B1(new_n607_), .B2(new_n386_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT42), .ZN(new_n634_));
  INV_X1    g433(.A(new_n386_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n591_), .A2(new_n449_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT99), .Z(G1327gat));
  INV_X1    g437(.A(new_n466_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n567_), .A2(new_n588_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n603_), .A2(new_n641_), .A3(new_n604_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n259_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n603_), .B2(new_n534_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n420_), .A2(KEYINPUT43), .A3(new_n535_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(KEYINPUT44), .A3(new_n646_), .A4(new_n640_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT43), .B1(new_n420_), .B2(new_n535_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n644_), .B(new_n534_), .C1(new_n404_), .C2(new_n419_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n654_), .B2(new_n641_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n649_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n608_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n643_), .B1(new_n657_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n642_), .A2(new_n659_), .A3(new_n410_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT45), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n649_), .A2(new_n410_), .A3(new_n655_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(G36gat), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n663_), .B(new_n666_), .ZN(G1329gat));
  XOR2_X1   g466(.A(KEYINPUT102), .B(G43gat), .Z(new_n668_));
  INV_X1    g467(.A(new_n642_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n403_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n416_), .A2(G43gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n656_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n642_), .B2(new_n635_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n656_), .A2(new_n386_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g475(.A(new_n567_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n587_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n606_), .A2(new_n639_), .A3(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT104), .B(G57gat), .Z(new_n680_));
  NOR3_X1   g479(.A1(new_n679_), .A2(new_n608_), .A3(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT105), .Z(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n537_), .A2(new_n678_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n608_), .B1(new_n685_), .B2(KEYINPUT103), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(KEYINPUT103), .B2(new_n685_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n683_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(new_n410_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G64gat), .B1(new_n679_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(G64gat), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT106), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n684_), .B2(new_n693_), .ZN(G1333gat));
  OAI21_X1  g493(.A(G71gat), .B1(new_n679_), .B2(new_n403_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT49), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n403_), .A2(G71gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n684_), .B2(new_n697_), .ZN(G1334gat));
  OAI21_X1  g497(.A(G78gat), .B1(new_n679_), .B2(new_n386_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT50), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n685_), .A2(new_n433_), .A3(new_n635_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT107), .ZN(G1335gat));
  NOR2_X1   g502(.A1(new_n603_), .A2(new_n604_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n677_), .A2(new_n587_), .A3(new_n639_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n259_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n653_), .A2(new_n705_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n259_), .A2(G85gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT108), .Z(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n710_), .B2(new_n712_), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n707_), .B2(new_n410_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n497_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n496_), .A2(G92gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n689_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n710_), .B2(new_n717_), .ZN(G1337gat));
  OAI21_X1  g517(.A(G99gat), .B1(new_n709_), .B2(new_n403_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n416_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n706_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g521(.A1(new_n653_), .A2(KEYINPUT109), .A3(new_n635_), .A4(new_n705_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n645_), .A2(new_n635_), .A3(new_n646_), .A4(new_n705_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n723_), .A2(new_n726_), .A3(KEYINPUT110), .A4(G106gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(KEYINPUT52), .A3(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n707_), .A2(new_n479_), .A3(new_n635_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n728_), .A3(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n731_), .A2(new_n737_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n547_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n550_), .A2(KEYINPUT55), .A3(new_n542_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT111), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n550_), .A2(new_n746_), .A3(KEYINPUT55), .A4(new_n542_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n559_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n750_));
  INV_X1    g549(.A(new_n560_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n574_), .A2(new_n575_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n580_), .B1(new_n753_), .B2(new_n569_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n568_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n581_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n757_), .A3(new_n559_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n750_), .A2(new_n751_), .A3(new_n756_), .A4(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n535_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n759_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(KEYINPUT113), .A3(new_n535_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n750_), .A2(new_n587_), .A3(new_n751_), .A4(new_n758_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n756_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n605_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n465_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n466_), .A2(new_n535_), .A3(new_n587_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n677_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n677_), .B2(new_n776_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n740_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n465_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n761_), .B2(new_n535_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n763_), .B(new_n534_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n765_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n771_), .B(KEYINPUT57), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n779_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT114), .A3(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n601_), .A2(new_n608_), .A3(new_n410_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n780_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n587_), .ZN(new_n791_));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n780_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n639_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n795_), .A2(new_n779_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n608_), .A2(new_n410_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n417_), .A4(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT115), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n802_), .A3(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n792_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n791_), .B1(new_n804_), .B2(new_n587_), .ZN(G1340gat));
  INV_X1    g604(.A(G120gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n677_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n790_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n806_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G120gat), .B1(new_n800_), .B2(new_n677_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1341gat));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n793_), .B2(new_n466_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT117), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n781_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g616(.A(G134gat), .B1(new_n790_), .B2(new_n605_), .ZN(new_n818_));
  INV_X1    g617(.A(G134gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n820_), .B2(new_n535_), .ZN(G1343gat));
  NAND4_X1  g620(.A1(new_n780_), .A2(new_n788_), .A3(new_n418_), .A4(new_n798_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n588_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT118), .B(G141gat), .Z(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1344gat));
  OR3_X1    g624(.A1(new_n822_), .A2(KEYINPUT120), .A3(new_n677_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n822_), .B2(new_n677_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT119), .B(G148gat), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1345gat));
  OR3_X1    g632(.A1(new_n822_), .A2(KEYINPUT121), .A3(new_n466_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT121), .B1(new_n822_), .B2(new_n466_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1346gat));
  NOR3_X1   g640(.A1(new_n822_), .A2(new_n203_), .A3(new_n534_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n780_), .A2(new_n788_), .A3(new_n418_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n605_), .A3(new_n798_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n203_), .B2(new_n844_), .ZN(G1347gat));
  NOR2_X1   g644(.A1(new_n689_), .A2(new_n259_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n417_), .B(new_n846_), .C1(new_n795_), .C2(new_n779_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n588_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n588_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(G169gat), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n285_), .A3(new_n587_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(G1348gat));
  NAND4_X1  g655(.A1(new_n780_), .A2(new_n788_), .A3(new_n417_), .A4(new_n846_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G176gat), .B1(new_n857_), .B2(new_n677_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n853_), .A2(new_n286_), .A3(new_n567_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT123), .ZN(G1349gat));
  NOR3_X1   g660(.A1(new_n847_), .A2(new_n781_), .A3(new_n293_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n857_), .A2(new_n466_), .ZN(new_n863_));
  INV_X1    g662(.A(G183gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n853_), .A2(new_n605_), .A3(new_n302_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n853_), .A2(new_n535_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT124), .B1(new_n867_), .B2(G190gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT124), .B(G190gat), .C1(new_n847_), .C2(new_n534_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT125), .B(new_n866_), .C1(new_n868_), .C2(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n843_), .A2(new_n846_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n588_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n677_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(G204gat), .Z(G1353gat));
  NAND2_X1  g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n465_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n883_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n876_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1354gat));
  NOR3_X1   g688(.A1(new_n876_), .A2(new_n468_), .A3(new_n534_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n843_), .A2(new_n605_), .A3(new_n846_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n468_), .B2(new_n891_), .ZN(G1355gat));
endmodule


