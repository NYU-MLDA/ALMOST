//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G85gat), .B(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(KEYINPUT9), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT6), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT65), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n203_), .A2(KEYINPUT8), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n221_), .B2(new_n212_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n212_), .B(KEYINPUT66), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n203_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G57gat), .B(G64gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G78gat), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n217_), .A2(new_n226_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n226_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n234_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n235_), .A2(new_n241_), .A3(KEYINPUT12), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT12), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n243_), .A3(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  AOI211_X1 g048(.A(new_n248_), .B(new_n249_), .C1(new_n242_), .C2(new_n244_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n235_), .A2(new_n241_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n249_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(G204gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT5), .B(G176gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n202_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT13), .A3(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G78gat), .B(G106gat), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G228gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n269_));
  AND3_X1   g068(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n269_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT89), .B(KEYINPUT1), .C1(new_n270_), .C2(new_n271_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  INV_X1    g078(.A(G141gat), .ZN(new_n280_));
  INV_X1    g079(.A(G148gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n281_), .A3(KEYINPUT3), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n279_), .A2(KEYINPUT90), .A3(KEYINPUT2), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT2), .B1(new_n279_), .B2(KEYINPUT90), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n287_), .B(KEYINPUT91), .C1(new_n288_), .C2(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n270_), .A2(new_n271_), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT92), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT92), .ZN(new_n298_));
  AOI211_X1 g097(.A(new_n298_), .B(new_n295_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n283_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT29), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(G197gat), .B(G204gat), .Z(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(KEYINPUT21), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT21), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT93), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n268_), .B1(new_n301_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n268_), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n310_), .B(new_n307_), .C1(new_n300_), .C2(KEYINPUT29), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n267_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n278_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n293_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n279_), .A2(KEYINPUT90), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n279_), .A2(KEYINPUT90), .A3(KEYINPUT2), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT91), .B1(new_n319_), .B2(new_n287_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n296_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n298_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n294_), .A2(KEYINPUT92), .A3(new_n296_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n313_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n308_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n310_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n301_), .A2(new_n268_), .A3(new_n308_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n266_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n312_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n325_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G22gat), .B(G50gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT28), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n331_), .B(new_n333_), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT94), .B1(new_n309_), .B2(new_n311_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n327_), .A2(new_n337_), .A3(new_n328_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .A4(new_n267_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(new_n329_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT96), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n338_), .A3(new_n267_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n334_), .B1(new_n343_), .B2(KEYINPUT95), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n335_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT97), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT97), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(new_n335_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G113gat), .ZN(new_n353_));
  INV_X1    g152(.A(G120gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n300_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT100), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n300_), .B(new_n355_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n356_), .B(new_n358_), .C1(new_n359_), .C2(new_n351_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n358_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G85gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n361_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  INV_X1    g171(.A(new_n306_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT23), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(KEYINPUT80), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(KEYINPUT23), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  INV_X1    g177(.A(G176gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT24), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT81), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(KEYINPUT24), .A3(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT78), .B(G190gat), .Z(new_n386_));
  INV_X1    g185(.A(KEYINPUT26), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n385_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT79), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(KEYINPUT79), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n383_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT82), .B1(new_n396_), .B2(G169gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G169gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n379_), .B(new_n397_), .C1(new_n398_), .C2(KEYINPUT82), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT83), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n376_), .A2(KEYINPUT23), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT84), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n401_), .B(KEYINPUT84), .C1(KEYINPUT23), .C2(new_n374_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n386_), .A2(G183gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n384_), .B(new_n400_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n373_), .B1(new_n395_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n398_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(G176gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n384_), .B1(new_n410_), .B2(KEYINPUT98), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n408_), .B(new_n411_), .C1(KEYINPUT98), .C2(new_n384_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n387_), .A2(G190gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n389_), .A2(new_n390_), .A3(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n402_), .A2(new_n403_), .A3(new_n385_), .A4(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n381_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n417_), .B2(new_n306_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n372_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n306_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n395_), .A2(new_n406_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT20), .B(new_n420_), .C1(new_n421_), .C2(new_n306_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n422_), .B2(new_n372_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT18), .B(G64gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(KEYINPUT32), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n372_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n432_));
  INV_X1    g231(.A(new_n427_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n370_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT101), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(new_n427_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n430_), .B(new_n433_), .C1(new_n422_), .C2(new_n429_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT99), .A3(new_n438_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n431_), .A2(KEYINPUT99), .A3(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n358_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n359_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n356_), .B1(new_n359_), .B2(new_n351_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n443_), .B(new_n366_), .C1(new_n444_), .C2(new_n358_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n369_), .A2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n369_), .A2(new_n446_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n441_), .A2(new_n445_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT101), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n370_), .A2(new_n450_), .A3(new_n428_), .A4(new_n434_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n436_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n348_), .A2(new_n350_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT102), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n348_), .A2(KEYINPUT102), .A3(new_n350_), .A4(new_n452_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT103), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n370_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n367_), .A2(KEYINPUT103), .A3(new_n369_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n439_), .A2(new_n440_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n423_), .A2(new_n433_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n437_), .A2(new_n463_), .A3(KEYINPUT27), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n344_), .A2(new_n329_), .A3(new_n340_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT96), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n349_), .B1(new_n470_), .B2(new_n335_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n350_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n460_), .B(new_n466_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n455_), .A2(new_n456_), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n421_), .B(KEYINPUT30), .Z(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT86), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT85), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G43gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n475_), .B2(KEYINPUT86), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n476_), .B(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n355_), .B(KEYINPUT31), .Z(new_n485_));
  AND2_X1   g284(.A1(new_n485_), .A2(KEYINPUT87), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n474_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n348_), .A2(new_n350_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT104), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n465_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n460_), .ZN(new_n492_));
  NOR4_X1   g291(.A1(new_n489_), .A2(new_n491_), .A3(new_n492_), .A4(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G15gat), .B(G22gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(G1gat), .A2(G8gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(KEYINPUT14), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT75), .ZN(new_n499_));
  XOR2_X1   g298(.A(G1gat), .B(G8gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  INV_X1    g302(.A(G43gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n501_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT77), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n501_), .B(new_n507_), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G229gat), .A3(G233gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(new_n378_), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(G197gat), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n515_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n495_), .A2(KEYINPUT105), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT105), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n493_), .B1(new_n474_), .B2(new_n487_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n525_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n265_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n234_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n501_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G183gat), .B(G211gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(KEYINPUT17), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n534_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n217_), .A2(new_n226_), .A3(new_n507_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n239_), .A2(new_n509_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(KEYINPUT35), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n545_), .A2(new_n546_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT69), .B(G134gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT36), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT71), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT71), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT70), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n550_), .A2(new_n553_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT37), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n567_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n562_), .A2(KEYINPUT74), .A3(new_n567_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n544_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n531_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G1gat), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n492_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n528_), .A2(new_n529_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n572_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n544_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n262_), .A2(new_n264_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n460_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n581_), .A2(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n583_), .A2(new_n589_), .A3(new_n590_), .ZN(G1324gat));
  INV_X1    g390(.A(G8gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n579_), .A2(new_n592_), .A3(new_n491_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n491_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G8gat), .B1(new_n588_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT39), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT39), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n588_), .B2(new_n487_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  INV_X1    g400(.A(G15gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n487_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n579_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(G1326gat));
  INV_X1    g404(.A(G22gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n579_), .A2(new_n606_), .A3(new_n489_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n489_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G22gat), .B1(new_n588_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(KEYINPUT42), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(KEYINPUT42), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT106), .Z(G1327gat));
  NOR2_X1   g412(.A1(new_n572_), .A2(new_n543_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n265_), .B(new_n615_), .C1(new_n526_), .C2(new_n530_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n460_), .A2(G29gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT110), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n587_), .A2(new_n544_), .A3(new_n525_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT107), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT43), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n570_), .A2(new_n577_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n495_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT43), .B1(new_n528_), .B2(new_n623_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n621_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT44), .ZN(new_n628_));
  INV_X1    g427(.A(new_n621_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n622_), .B1(new_n495_), .B2(new_n624_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n528_), .A2(KEYINPUT43), .A3(new_n623_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT44), .B(new_n629_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT108), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT108), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n634_), .A3(KEYINPUT44), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n628_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n492_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n637_), .A2(KEYINPUT109), .A3(G29gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT109), .B1(new_n637_), .B2(G29gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n619_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  OAI21_X1  g439(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n594_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n632_), .A2(KEYINPUT108), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n634_), .B1(new_n627_), .B2(KEYINPUT44), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n531_), .A2(new_n648_), .A3(new_n491_), .A4(new_n614_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n616_), .A2(KEYINPUT45), .A3(new_n648_), .A4(new_n491_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n647_), .A2(new_n653_), .A3(KEYINPUT111), .A4(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT111), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n654_), .A2(KEYINPUT111), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n633_), .A2(new_n635_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n648_), .B1(new_n658_), .B2(new_n643_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(new_n652_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n656_), .B(new_n657_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n655_), .A2(new_n661_), .ZN(G1329gat));
  NAND3_X1  g461(.A1(new_n636_), .A2(G43gat), .A3(new_n603_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n616_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n504_), .B1(new_n664_), .B2(new_n487_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT47), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1330gat));
  NAND2_X1  g469(.A1(new_n489_), .A2(new_n506_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT112), .Z(new_n672_));
  NOR2_X1   g471(.A1(new_n664_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT113), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n636_), .A2(new_n489_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n674_), .B(new_n675_), .C1(new_n676_), .C2(new_n506_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n506_), .B1(new_n636_), .B2(new_n489_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT113), .B1(new_n678_), .B2(new_n673_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1331gat));
  NAND4_X1  g479(.A1(new_n495_), .A2(new_n586_), .A3(new_n265_), .A4(new_n529_), .ZN(new_n681_));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n460_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n528_), .A2(new_n525_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT114), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n265_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n578_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n492_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n683_), .B1(new_n688_), .B2(new_n682_), .ZN(G1332gat));
  INV_X1    g488(.A(G64gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n690_), .A3(new_n491_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G64gat), .B1(new_n681_), .B2(new_n594_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT48), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n695_), .A3(new_n603_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G71gat), .B1(new_n681_), .B2(new_n487_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT49), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1334gat));
  INV_X1    g498(.A(G78gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(new_n700_), .A3(new_n489_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G78gat), .B1(new_n681_), .B2(new_n608_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1335gat));
  NAND3_X1  g503(.A1(new_n265_), .A2(new_n544_), .A3(new_n529_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT115), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n460_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n686_), .A2(new_n614_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n492_), .A2(new_n205_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT116), .ZN(G1336gat));
  NOR3_X1   g512(.A1(new_n708_), .A2(new_n206_), .A3(new_n594_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n686_), .A2(new_n491_), .A3(new_n614_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n206_), .ZN(G1337gat));
  NAND2_X1  g515(.A1(new_n603_), .A2(new_n214_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n707_), .A2(new_n603_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT117), .A3(G99gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT117), .B1(new_n718_), .B2(G99gat), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n710_), .A2(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  INV_X1    g522(.A(new_n706_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n489_), .B(new_n724_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT118), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n723_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(G106gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT118), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(KEYINPUT52), .A3(new_n727_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n686_), .A2(new_n213_), .A3(new_n489_), .A4(new_n614_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n730_), .A2(new_n733_), .A3(new_n734_), .A4(new_n736_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1339gat));
  INV_X1    g539(.A(KEYINPUT120), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n623_), .A2(new_n543_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n262_), .A2(new_n264_), .A3(new_n529_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n587_), .A2(KEYINPUT120), .A3(new_n529_), .A4(new_n578_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT54), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n741_), .B(new_n747_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n242_), .A2(new_n249_), .A3(new_n244_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n245_), .A2(KEYINPUT55), .A3(new_n246_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n258_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT121), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n755_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n516_), .A2(new_n512_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n511_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(new_n521_), .C1(new_n763_), .C2(new_n512_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n524_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n755_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n260_), .B1(new_n767_), .B2(KEYINPUT121), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n761_), .A2(new_n768_), .A3(KEYINPUT58), .A4(new_n766_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n624_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n263_), .B2(new_n259_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n758_), .A2(new_n760_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n525_), .A2(new_n259_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n778_), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n572_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n572_), .C1(new_n780_), .C2(new_n774_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n572_), .B1(new_n780_), .B2(new_n774_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n773_), .A2(new_n779_), .A3(new_n783_), .A4(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n749_), .B1(new_n787_), .B2(new_n544_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n608_), .A2(new_n603_), .A3(new_n594_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n460_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n525_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n790_), .B(KEYINPUT59), .Z(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(new_n529_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g593(.A(G120gat), .B1(new_n792_), .B2(new_n587_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n354_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n790_), .B(new_n796_), .C1(KEYINPUT60), .C2(new_n354_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n790_), .B2(new_n543_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT123), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n792_), .A2(new_n544_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g601(.A(G134gat), .B1(new_n790_), .B2(new_n585_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n792_), .A2(new_n623_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n787_), .A2(new_n544_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n749_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n608_), .A2(new_n603_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n492_), .A3(new_n594_), .A4(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT124), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n809_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n788_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT124), .A3(new_n492_), .A4(new_n594_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n525_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n265_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n543_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  INV_X1    g622(.A(G162gat), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n824_), .B(new_n623_), .C1(new_n812_), .C2(new_n815_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n816_), .A2(new_n585_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n824_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n572_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT125), .B1(new_n829_), .B2(G162gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n828_), .B2(new_n830_), .ZN(G1347gat));
  NOR3_X1   g630(.A1(new_n788_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n594_), .A2(new_n492_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n529_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n835_), .B2(new_n378_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n837_), .B(new_n839_), .C1(new_n409_), .C2(new_n836_), .ZN(G1348gat));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n587_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n379_), .ZN(G1349gat));
  NOR2_X1   g641(.A1(new_n834_), .A2(new_n544_), .ZN(new_n843_));
  MUX2_X1   g642(.A(G183gat), .B(new_n389_), .S(new_n843_), .Z(G1350gat));
  OAI21_X1  g643(.A(G190gat), .B1(new_n834_), .B2(new_n623_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n585_), .A2(new_n390_), .A3(new_n413_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n834_), .B2(new_n846_), .ZN(G1351gat));
  NAND2_X1  g646(.A1(new_n814_), .A2(new_n833_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n525_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g650(.A1(new_n848_), .A2(new_n587_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n853_));
  AND2_X1   g652(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n852_), .B2(new_n853_), .ZN(G1353gat));
  NAND2_X1  g655(.A1(new_n849_), .A2(new_n543_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n857_), .B2(new_n858_), .ZN(G1354gat));
  NAND3_X1  g660(.A1(new_n849_), .A2(G218gat), .A3(new_n624_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n848_), .A2(new_n572_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(G218gat), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT127), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n862_), .B(KEYINPUT127), .C1(G218gat), .C2(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1355gat));
endmodule


