//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT66), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT7), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(KEYINPUT67), .A3(new_n216_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT8), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n207_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n216_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n213_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT65), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(KEYINPUT65), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n231_), .B(new_n232_), .C1(new_n227_), .C2(new_n213_), .ZN(new_n233_));
  OAI221_X1 g032(.A(new_n207_), .B1(G106gat), .B2(new_n226_), .C1(new_n233_), .C2(new_n215_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n225_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n225_), .B2(new_n234_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  OAI22_X1  g042(.A1(new_n241_), .A2(new_n242_), .B1(new_n243_), .B2(KEYINPUT12), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n245_));
  AND2_X1   g044(.A1(new_n225_), .A2(new_n234_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(new_n240_), .ZN(new_n247_));
  INV_X1    g046(.A(G230gat), .ZN(new_n248_));
  INV_X1    g047(.A(G233gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n244_), .B(new_n247_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n249_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G176gat), .B(G204gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G120gat), .B(G148gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n253_), .A2(new_n258_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT76), .B(G22gat), .ZN(new_n268_));
  INV_X1    g067(.A(G15gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT77), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G29gat), .B(G36gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G43gat), .B(G50gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT15), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n277_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G229gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n279_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n285_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G169gat), .B(G197gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n297_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n267_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT31), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT23), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(G183gat), .A3(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G183gat), .ZN(new_n312_));
  INV_X1    g111(.A(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  AND2_X1   g116(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT26), .B1(new_n313_), .B2(KEYINPUT80), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(G190gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n308_), .A2(new_n310_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT24), .A3(new_n316_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n321_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT30), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G43gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT81), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(new_n269_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G71gat), .B(G99gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n336_), .B(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n306_), .B1(new_n342_), .B2(KEYINPUT82), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(KEYINPUT82), .B2(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n342_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n306_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n305_), .ZN(new_n349_));
  AND2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350_));
  INV_X1    g149(.A(G141gat), .ZN(new_n351_));
  INV_X1    g150(.A(G148gat), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n350_), .A2(KEYINPUT1), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G155gat), .B(G162gat), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n353_), .B(new_n354_), .C1(KEYINPUT1), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n350_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n349_), .B1(new_n367_), .B2(KEYINPUT95), .ZN(new_n368_));
  INV_X1    g167(.A(new_n354_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n371_), .A2(new_n353_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n305_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n374_), .A3(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(new_n372_), .A2(new_n305_), .A3(KEYINPUT4), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n368_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT0), .B(G57gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n387_), .A3(new_n380_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n367_), .B2(KEYINPUT29), .ZN(new_n391_));
  INV_X1    g190(.A(G197gat), .ZN(new_n392_));
  AND2_X1   g191(.A1(KEYINPUT83), .A2(G204gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(KEYINPUT83), .A2(G204gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G197gat), .A2(G204gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT21), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(G197gat), .B1(new_n393_), .B2(new_n394_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT21), .ZN(new_n399_));
  INV_X1    g198(.A(G204gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(G197gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G211gat), .ZN(new_n404_));
  INV_X1    g203(.A(G218gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G211gat), .A2(G218gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n397_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT83), .B(G204gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n401_), .B1(new_n411_), .B2(G197gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n407_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n398_), .A2(new_n402_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n413_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT84), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n391_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT85), .B1(new_n372_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n367_), .A2(new_n423_), .A3(KEYINPUT29), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n390_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(KEYINPUT86), .A3(new_n390_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n420_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G78gat), .B(G106gat), .Z(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT87), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT88), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(KEYINPUT89), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n372_), .A2(new_n421_), .ZN(new_n435_));
  INV_X1    g234(.A(G50gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT28), .B(G22gat), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n438_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n425_), .A2(KEYINPUT86), .A3(new_n390_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT86), .B1(new_n425_), .B2(new_n390_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n433_), .B(new_n419_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n434_), .B(new_n442_), .C1(new_n444_), .C2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n419_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n432_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n451_), .A2(KEYINPUT90), .A3(new_n447_), .A4(new_n441_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n449_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G92gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT18), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT26), .B(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n322_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n320_), .A2(KEYINPUT92), .A3(new_n316_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT92), .B1(new_n320_), .B2(new_n316_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n311_), .A2(KEYINPUT93), .A3(new_n314_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT93), .B1(new_n311_), .B2(new_n314_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n470_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n409_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n466_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n418_), .A2(new_n334_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n465_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n414_), .A2(new_n417_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n473_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n477_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n475_), .A4(new_n471_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n484_), .A2(new_n409_), .B1(new_n487_), .B2(new_n469_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n334_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n464_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n461_), .B1(new_n483_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n469_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n482_), .B(KEYINPUT20), .C1(new_n492_), .C2(new_n418_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n464_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n418_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n418_), .A2(new_n334_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT20), .A4(new_n465_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n460_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(KEYINPUT94), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT27), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n497_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n461_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n464_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n488_), .A2(new_n489_), .A3(new_n465_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n460_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n491_), .A2(new_n507_), .A3(KEYINPUT27), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n491_), .A2(new_n507_), .A3(KEYINPUT99), .A4(KEYINPUT27), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NOR4_X1   g311(.A1(new_n348_), .A2(new_n389_), .A3(new_n456_), .A4(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n504_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n389_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n456_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT100), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n456_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n505_), .A2(new_n506_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n461_), .A2(KEYINPUT32), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n522_), .B(new_n515_), .C1(new_n521_), .C2(new_n501_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n379_), .A2(KEYINPUT33), .A3(new_n387_), .A4(new_n380_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(KEYINPUT96), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(KEYINPUT96), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n368_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n385_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT98), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n531_), .A3(new_n385_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n525_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n388_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n499_), .A2(new_n503_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n519_), .B1(new_n523_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n514_), .A2(new_n456_), .A3(KEYINPUT100), .A4(new_n515_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n518_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n513_), .B1(new_n541_), .B2(new_n348_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  INV_X1    g342(.A(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT73), .B(G134gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n246_), .B2(new_n282_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n225_), .A2(new_n234_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n283_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n551_), .A2(new_n556_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n558_), .B2(new_n289_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n555_), .B(new_n554_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n549_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT75), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n571_), .B(new_n549_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n240_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n279_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G211gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT16), .B(G183gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT17), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT78), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n578_), .A2(new_n586_), .A3(new_n582_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(KEYINPUT78), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT79), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n575_), .A2(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n302_), .A2(new_n542_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR4_X1   g394(.A1(new_n302_), .A2(new_n542_), .A3(new_n592_), .A4(KEYINPUT101), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(G1gat), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n598_), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n389_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n593_), .A2(new_n594_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n271_), .B(new_n389_), .C1(new_n601_), .C2(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n589_), .ZN(new_n606_));
  NOR4_X1   g405(.A1(new_n302_), .A2(new_n542_), .A3(new_n568_), .A4(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT103), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n389_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G1gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n602_), .A2(KEYINPUT104), .A3(new_n603_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT104), .B1(new_n602_), .B2(new_n603_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n202_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(KEYINPUT105), .A3(new_n605_), .A4(new_n610_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1324gat));
  AOI21_X1  g417(.A(new_n272_), .B1(new_n607_), .B2(new_n512_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n272_), .B(new_n512_), .C1(new_n601_), .C2(new_n596_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g423(.A(new_n348_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n593_), .A2(new_n269_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n269_), .B1(new_n608_), .B2(new_n625_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n608_), .B2(new_n456_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT42), .Z(new_n634_));
  NAND3_X1  g433(.A1(new_n593_), .A2(new_n632_), .A3(new_n456_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1327gat));
  NAND2_X1  g435(.A1(new_n541_), .A2(new_n348_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n513_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  INV_X1    g439(.A(new_n575_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT43), .B1(new_n542_), .B2(new_n575_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n302_), .A2(new_n591_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n389_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n640_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n542_), .A2(KEYINPUT43), .A3(new_n575_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n644_), .A2(KEYINPUT108), .A3(new_n645_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n652_), .A2(KEYINPUT110), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n647_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(G29gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n568_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n542_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n645_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n389_), .A2(new_n660_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT111), .ZN(new_n666_));
  OAI22_X1  g465(.A1(new_n659_), .A2(new_n660_), .B1(new_n664_), .B2(new_n666_), .ZN(G1328gat));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n668_), .A3(new_n512_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n646_), .A2(new_n512_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n672_), .B2(new_n668_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT46), .B(new_n670_), .C1(new_n672_), .C2(new_n668_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND2_X1  g476(.A1(new_n646_), .A2(G43gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n348_), .B(new_n678_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G43gat), .B1(new_n663_), .B2(new_n625_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT47), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n625_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(new_n680_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n681_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n663_), .B2(new_n456_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n436_), .B(new_n519_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n646_), .ZN(G1331gat));
  NOR2_X1   g489(.A1(new_n542_), .A2(new_n301_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n591_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n267_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n693_), .A3(new_n661_), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n515_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n691_), .A2(new_n693_), .A3(new_n575_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(new_n515_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n695_), .B2(new_n698_), .ZN(G1332gat));
  OAI21_X1  g498(.A(G64gat), .B1(new_n694_), .B2(new_n514_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT48), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n514_), .A2(G64gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n697_), .B2(new_n702_), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n694_), .B2(new_n348_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT49), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n697_), .A2(G71gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n348_), .B2(new_n706_), .ZN(G1334gat));
  OAI21_X1  g506(.A(G78gat), .B1(new_n694_), .B2(new_n519_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT50), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n519_), .A2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n697_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT112), .ZN(G1335gat));
  INV_X1    g511(.A(G85gat), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n267_), .A2(new_n301_), .A3(new_n591_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n662_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n715_), .B2(new_n515_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT113), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n644_), .A2(new_n714_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(new_n713_), .A3(new_n515_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1336gat));
  INV_X1    g519(.A(G92gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n715_), .B2(new_n514_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT114), .Z(new_n723_));
  INV_X1    g522(.A(new_n718_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n514_), .A2(new_n721_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n718_), .B2(new_n348_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n348_), .A2(new_n226_), .ZN(new_n729_));
  OAI221_X1 g528(.A(new_n727_), .B1(KEYINPUT115), .B2(new_n728_), .C1(new_n715_), .C2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(KEYINPUT115), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1338gat));
  OR3_X1    g531(.A1(new_n715_), .A2(G106gat), .A3(new_n519_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n724_), .A2(new_n456_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G106gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G106gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g538(.A1(new_n267_), .A2(new_n575_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n591_), .A2(new_n300_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT116), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n740_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n259_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n250_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n244_), .A2(KEYINPUT55), .A3(new_n247_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n251_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n251_), .A2(new_n751_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n244_), .A2(KEYINPUT55), .A3(new_n247_), .A4(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n749_), .A2(new_n752_), .A3(KEYINPUT118), .A4(new_n754_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n258_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n747_), .B1(new_n759_), .B2(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n286_), .A2(new_n292_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n291_), .A2(new_n287_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n297_), .A3(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT120), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n298_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n757_), .A2(new_n766_), .A3(new_n258_), .A4(new_n758_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n760_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n760_), .A2(KEYINPUT58), .A3(new_n765_), .A4(new_n767_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n641_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n259_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n759_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n757_), .A2(new_n258_), .A3(new_n774_), .A4(new_n758_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n301_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n261_), .A2(new_n765_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n773_), .B1(new_n780_), .B2(new_n661_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT57), .B(new_n568_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n772_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n746_), .B1(new_n783_), .B2(new_n606_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n456_), .A2(new_n512_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n625_), .A2(new_n389_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G113gat), .B1(new_n787_), .B2(new_n301_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n787_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n300_), .B1(new_n759_), .B2(new_n775_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n790_), .A2(new_n777_), .B1(new_n261_), .B2(new_n765_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT57), .B1(new_n791_), .B2(new_n568_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n780_), .A2(new_n773_), .A3(new_n661_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n591_), .B1(new_n794_), .B2(new_n772_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n795_), .A2(new_n746_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n789_), .A2(KEYINPUT59), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n301_), .A2(G113gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n788_), .B1(new_n798_), .B2(new_n799_), .ZN(G1340gat));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n797_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n267_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n802_), .C1(new_n803_), .C2(new_n787_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT121), .B(G120gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n267_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n787_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n807_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g609(.A(G127gat), .B1(new_n787_), .B2(new_n591_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n589_), .A2(G127gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n798_), .B2(new_n812_), .ZN(G1342gat));
  AOI21_X1  g612(.A(G134gat), .B1(new_n787_), .B2(new_n568_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n641_), .A2(G134gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n798_), .B2(new_n815_), .ZN(G1343gat));
  NOR3_X1   g615(.A1(new_n625_), .A2(new_n519_), .A3(new_n512_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n589_), .B1(new_n794_), .B2(new_n772_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n389_), .B(new_n817_), .C1(new_n818_), .C2(new_n746_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n300_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(new_n351_), .ZN(G1344gat));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n267_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(new_n352_), .ZN(G1345gat));
  OAI21_X1  g622(.A(KEYINPUT122), .B1(new_n819_), .B2(new_n692_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n783_), .A2(new_n606_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n746_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n515_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n591_), .A4(new_n817_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n824_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1346gat));
  NOR3_X1   g632(.A1(new_n819_), .A2(new_n544_), .A3(new_n575_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n827_), .A2(new_n568_), .A3(new_n817_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n544_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n348_), .A2(new_n389_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n519_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n512_), .B(new_n839_), .C1(new_n795_), .C2(new_n746_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G169gat), .B1(new_n840_), .B2(new_n300_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n300_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n319_), .B2(new_n318_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .ZN(G1348gat));
  OAI21_X1  g646(.A(new_n317_), .B1(new_n840_), .B2(new_n267_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT124), .B(new_n317_), .C1(new_n840_), .C2(new_n267_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n784_), .A2(new_n514_), .A3(new_n838_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n267_), .A2(new_n317_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n850_), .A2(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  NOR3_X1   g653(.A1(new_n840_), .A2(new_n322_), .A3(new_n606_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n591_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n312_), .ZN(G1350gat));
  OAI21_X1  g656(.A(G190gat), .B1(new_n840_), .B2(new_n575_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n568_), .A2(new_n467_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n796_), .A2(new_n512_), .A3(new_n839_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n858_), .A2(new_n861_), .A3(KEYINPUT125), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1351gat));
  NAND2_X1  g665(.A1(new_n825_), .A2(new_n826_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n625_), .A2(new_n389_), .A3(new_n519_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(KEYINPUT126), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(KEYINPUT126), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n867_), .A2(new_n512_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n300_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n392_), .ZN(G1352gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n267_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n411_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n400_), .B2(new_n876_), .ZN(G1353gat));
  AOI21_X1  g677(.A(new_n514_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(new_n589_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT63), .B(G211gat), .Z(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT127), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n884_), .A3(new_n404_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n872_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n784_), .A2(new_n514_), .A3(new_n870_), .A4(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(new_n589_), .A4(new_n881_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n883_), .A2(new_n885_), .A3(new_n889_), .ZN(G1354gat));
  AOI21_X1  g689(.A(G218gat), .B1(new_n887_), .B2(new_n568_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n873_), .A2(new_n405_), .A3(new_n575_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1355gat));
endmodule


