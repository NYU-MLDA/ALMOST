//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n205_), .B(new_n206_), .C1(G183gat), .C2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n212_), .B2(KEYINPUT22), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n207_), .B(new_n208_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT81), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n203_), .B(KEYINPUT23), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT80), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n222_), .A2(new_n223_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n216_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT87), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n231_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n209_), .A2(new_n214_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n217_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n223_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n226_), .A3(new_n219_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n239_), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT20), .B(new_n240_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT19), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n231_), .B2(new_n239_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n255_), .A2(new_n257_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G8gat), .B(G36gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  AOI21_X1  g067(.A(new_n202_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n254_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n261_), .B1(new_n270_), .B2(new_n260_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT20), .B1(new_n231_), .B2(new_n239_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n249_), .B(new_n250_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n242_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n274_), .B2(new_n239_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n275_), .B2(new_n261_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n268_), .B(KEYINPUT95), .Z(new_n277_));
  NOR3_X1   g076(.A1(new_n276_), .A2(KEYINPUT96), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279_));
  INV_X1    g078(.A(new_n271_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n277_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n269_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G228gat), .A2(G233gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT88), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n239_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G141gat), .ZN(new_n290_));
  INV_X1    g089(.A(G148gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n289_), .A2(KEYINPUT2), .B1(new_n292_), .B2(KEYINPUT3), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n288_), .B(new_n294_), .ZN(new_n295_));
  OAI221_X1 g094(.A(new_n293_), .B1(KEYINPUT3), .B2(new_n292_), .C1(new_n295_), .C2(KEYINPUT2), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT86), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(KEYINPUT1), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n295_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n292_), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n239_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n287_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n287_), .A2(new_n307_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT90), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n314_), .A3(new_n311_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n305_), .A2(new_n316_), .A3(new_n306_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n300_), .A2(new_n304_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT28), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n311_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n308_), .A2(new_n309_), .A3(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n313_), .A2(new_n315_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n312_), .A2(KEYINPUT89), .A3(new_n328_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n308_), .A2(new_n331_), .A3(new_n309_), .A4(new_n327_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(new_n325_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341_));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n305_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(KEYINPUT84), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(new_n343_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n318_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n305_), .A2(new_n348_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(KEYINPUT4), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n355_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n340_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n340_), .A3(new_n358_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n258_), .A2(new_n262_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n268_), .C1(new_n275_), .C2(new_n261_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n255_), .A2(new_n257_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n268_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n202_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n284_), .A2(new_n335_), .A3(new_n363_), .A4(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n364_), .B1(new_n275_), .B2(new_n261_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n268_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n359_), .A2(KEYINPUT33), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n373_), .A2(new_n365_), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n340_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n353_), .A2(KEYINPUT4), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(KEYINPUT4), .B2(new_n351_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT94), .B1(new_n378_), .B2(new_n356_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n352_), .A2(new_n354_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n355_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n376_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n360_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n268_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n263_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n360_), .A2(new_n361_), .B1(new_n281_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n375_), .A2(new_n385_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n370_), .B1(new_n390_), .B2(new_n335_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n231_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n348_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n394_), .A2(new_n349_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n396_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n396_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT27), .B1(new_n373_), .B2(new_n365_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT96), .B1(new_n276_), .B2(new_n277_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n281_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n409_), .B2(new_n269_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n315_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n412_), .A2(new_n313_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n405_), .A2(new_n362_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n284_), .A2(new_n413_), .A3(new_n414_), .A4(new_n369_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT97), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n391_), .A2(new_n405_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G141gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G169gat), .B(G197gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  XNOR2_X1  g220(.A(G29gat), .B(G36gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT74), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n423_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT15), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G15gat), .B(G22gat), .ZN(new_n429_));
  INV_X1    g228(.A(G1gat), .ZN(new_n430_));
  INV_X1    g229(.A(G8gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT14), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G8gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n426_), .A2(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G229gat), .A2(G233gat), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n426_), .B(new_n435_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n421_), .B1(new_n444_), .B2(KEYINPUT79), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446_));
  INV_X1    g245(.A(new_n421_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n443_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n450_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(KEYINPUT65), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT67), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n455_), .A2(new_n465_), .A3(new_n459_), .A4(new_n462_), .ZN(new_n466_));
  INV_X1    g265(.A(G85gat), .ZN(new_n467_));
  INV_X1    g266(.A(G92gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(KEYINPUT8), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n466_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n459_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT8), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT64), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n478_), .A2(new_n483_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n469_), .A2(KEYINPUT9), .A3(new_n470_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n455_), .A2(new_n462_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT66), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n455_), .A2(new_n462_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n484_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n487_), .A2(new_n486_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n477_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT69), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G71gat), .A2(G78gat), .ZN(new_n500_));
  INV_X1    g299(.A(G71gat), .ZN(new_n501_));
  INV_X1    g300(.A(G78gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n500_), .B(new_n503_), .C1(new_n497_), .C2(KEYINPUT11), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n499_), .B(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n496_), .A2(KEYINPUT12), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n477_), .A2(KEYINPUT68), .A3(new_n495_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT68), .B1(new_n477_), .B2(new_n495_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n489_), .A2(new_n494_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n472_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n463_), .B2(KEYINPUT67), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n516_), .A2(new_n466_), .B1(new_n475_), .B2(KEYINPUT8), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n505_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n477_), .A2(KEYINPUT68), .A3(new_n495_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n512_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n522_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n521_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G120gat), .B(G148gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n533_), .B(KEYINPUT71), .Z(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT72), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n524_), .A2(new_n528_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n534_), .C1(new_n540_), .C2(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n418_), .A2(new_n449_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT73), .Z(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT75), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n508_), .A2(new_n509_), .A3(new_n426_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n428_), .B2(new_n496_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(KEYINPUT75), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n552_), .A2(KEYINPUT75), .A3(new_n550_), .A4(new_n554_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT36), .Z(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n564_), .A2(new_n567_), .A3(KEYINPUT37), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n564_), .B2(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n435_), .B(KEYINPUT76), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n505_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n574_), .B1(new_n578_), .B2(KEYINPUT17), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n574_), .A2(KEYINPUT17), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT77), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n581_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n570_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT78), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n546_), .A2(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n588_), .A2(G1gat), .A3(new_n363_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n564_), .A2(new_n567_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n418_), .A2(new_n584_), .A3(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n545_), .A2(new_n449_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n363_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n592_), .A3(new_n597_), .ZN(G1324gat));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n594_), .A2(new_n595_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n410_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n602_), .B2(G8gat), .ZN(new_n603_));
  AOI211_X1 g402(.A(KEYINPUT39), .B(new_n431_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n431_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n603_), .A2(new_n604_), .B1(new_n588_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n596_), .B2(new_n405_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n611_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n405_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n398_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n612_), .B(new_n613_), .C1(new_n588_), .C2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g416(.A(G22gat), .B1(new_n596_), .B2(new_n413_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT42), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(KEYINPUT42), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n413_), .A2(G22gat), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n619_), .A2(new_n620_), .B1(new_n588_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT102), .Z(G1327gat));
  INV_X1    g422(.A(new_n593_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n585_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n546_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n362_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n570_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n391_), .A2(new_n405_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n415_), .A2(new_n417_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  INV_X1    g432(.A(new_n570_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n545_), .A2(new_n449_), .A3(new_n585_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n636_), .A2(KEYINPUT103), .A3(KEYINPUT44), .A4(new_n637_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n637_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n640_), .A2(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n362_), .A2(G29gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n628_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  INV_X1    g445(.A(KEYINPUT46), .ZN(new_n647_));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n644_), .B2(new_n601_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n410_), .A2(KEYINPUT104), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n410_), .A2(KEYINPUT104), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n627_), .A2(new_n648_), .A3(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT45), .Z(new_n654_));
  OAI21_X1  g453(.A(new_n647_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n640_), .A2(new_n641_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n643_), .A2(new_n642_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G36gat), .B1(new_n658_), .B2(new_n410_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n653_), .B(KEYINPUT45), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(KEYINPUT46), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n661_), .ZN(G1329gat));
  INV_X1    g461(.A(G43gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n626_), .B2(new_n405_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n614_), .A2(G43gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n658_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT47), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n664_), .C1(new_n658_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1330gat));
  OR3_X1    g469(.A1(new_n626_), .A2(G50gat), .A3(new_n413_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n644_), .A2(KEYINPUT105), .A3(new_n335_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G50gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT105), .B1(new_n644_), .B2(new_n335_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1331gat));
  AND3_X1   g474(.A1(new_n594_), .A2(new_n449_), .A3(new_n545_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(G57gat), .A3(new_n362_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT106), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT106), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n445_), .A2(new_n448_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n418_), .A2(new_n680_), .A3(new_n544_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n587_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n362_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n678_), .A2(new_n679_), .A3(new_n684_), .ZN(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n676_), .B2(new_n652_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n652_), .A2(new_n686_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(new_n692_));
  OAI22_X1  g491(.A1(new_n689_), .A2(new_n690_), .B1(new_n682_), .B2(new_n692_), .ZN(G1333gat));
  NAND3_X1  g492(.A1(new_n683_), .A2(new_n501_), .A3(new_n614_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n501_), .B1(new_n676_), .B2(new_n614_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1334gat));
  NAND3_X1  g498(.A1(new_n683_), .A2(new_n502_), .A3(new_n335_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n502_), .B1(new_n676_), .B2(new_n335_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT50), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT50), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1335gat));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n629_), .A2(new_n635_), .A3(new_n706_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n544_), .A2(new_n680_), .A3(new_n585_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT109), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n636_), .A2(KEYINPUT108), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n708_), .A4(new_n707_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n362_), .A2(G85gat), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT110), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n681_), .A2(new_n625_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n467_), .B1(new_n718_), .B2(new_n363_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1336gat));
  INV_X1    g521(.A(new_n718_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n468_), .A3(new_n601_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n711_), .A2(new_n652_), .A3(new_n714_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n468_), .ZN(G1337gat));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n614_), .A3(new_n714_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G99gat), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n723_), .A2(new_n614_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n636_), .A2(new_n335_), .A3(new_n708_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT52), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n718_), .A2(G106gat), .A3(new_n413_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT112), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n737_), .A2(new_n739_), .A3(new_n743_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  NAND2_X1  g544(.A1(new_n680_), .A2(new_n534_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n521_), .B(new_n506_), .C1(new_n527_), .C2(KEYINPUT12), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n525_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n506_), .B1(new_n527_), .B2(KEYINPUT12), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n521_), .A2(new_n522_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(KEYINPUT55), .A3(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n512_), .B2(new_n523_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n748_), .B(new_n750_), .C1(new_n753_), .C2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n536_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT55), .B1(new_n751_), .B2(new_n752_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n512_), .A2(new_n523_), .A3(new_n754_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n748_), .B1(new_n762_), .B2(new_n750_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n758_), .A2(new_n759_), .A3(new_n763_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n760_), .A2(new_n761_), .B1(new_n525_), .B2(new_n749_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n536_), .B1(new_n765_), .B2(new_n748_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n750_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT113), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n747_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n440_), .A2(new_n438_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n447_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n538_), .A2(new_n541_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n593_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n534_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n759_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n757_), .A4(new_n756_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n570_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n777_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n781_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n776_), .A2(KEYINPUT57), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n776_), .B2(KEYINPUT57), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n746_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n775_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n624_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT114), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n787_), .A2(new_n789_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n584_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n680_), .B(new_n584_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n544_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n797_), .B2(new_n544_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n796_), .A2(new_n803_), .ZN(new_n804_));
  NOR4_X1   g603(.A1(new_n601_), .A2(new_n363_), .A3(new_n335_), .A4(new_n405_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n680_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT57), .B(new_n624_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n784_), .B(new_n782_), .C1(new_n764_), .C2(new_n769_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n634_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n780_), .A2(new_n782_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n776_), .A2(KEYINPUT57), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n584_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n802_), .B1(new_n815_), .B2(KEYINPUT116), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(KEYINPUT116), .B2(new_n815_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n805_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(G113gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n680_), .A2(KEYINPUT117), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(G113gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n808_), .B1(new_n822_), .B2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n821_), .B2(new_n544_), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n832_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT119), .B1(new_n807_), .B2(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n835_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(new_n836_), .B2(new_n837_), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n821_), .B2(new_n584_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n584_), .A2(G127gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n806_), .B2(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n821_), .B2(new_n570_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n624_), .A2(G134gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n806_), .B2(new_n843_), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n802_), .B1(new_n795_), .B2(new_n584_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n614_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n652_), .A2(new_n363_), .A3(new_n413_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n680_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT120), .B(G141gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n545_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n585_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  INV_X1    g655(.A(G162gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n857_), .A3(new_n593_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n848_), .A2(new_n634_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n857_), .ZN(G1347gat));
  NAND2_X1  g659(.A1(new_n652_), .A2(new_n414_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n861_), .A2(new_n335_), .A3(new_n449_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n817_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G169gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n817_), .A2(new_n209_), .A3(new_n862_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n864_), .A2(KEYINPUT121), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n212_), .B1(new_n817_), .B2(new_n862_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT62), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n866_), .B(new_n867_), .C1(new_n868_), .C2(new_n871_), .ZN(G1348gat));
  OAI21_X1  g671(.A(KEYINPUT122), .B1(new_n845_), .B2(new_n335_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT114), .B1(new_n792_), .B2(new_n793_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n813_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n585_), .B1(new_n876_), .B2(new_n794_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n874_), .B(new_n413_), .C1(new_n877_), .C2(new_n802_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n861_), .A2(new_n544_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n214_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n861_), .A2(new_n335_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n817_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n545_), .A2(new_n214_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT123), .B1(new_n881_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  INV_X1    g686(.A(new_n880_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n873_), .B2(new_n878_), .ZN(new_n889_));
  OAI221_X1 g688(.A(new_n887_), .B1(new_n883_), .B2(new_n884_), .C1(new_n889_), .C2(new_n214_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n890_), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n883_), .A2(new_n224_), .A3(new_n584_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n879_), .A2(new_n414_), .A3(new_n585_), .A4(new_n652_), .ZN(new_n893_));
  INV_X1    g692(.A(G183gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n883_), .B2(new_n570_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n593_), .A2(new_n225_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n883_), .B2(new_n897_), .ZN(G1351gat));
  XOR2_X1   g697(.A(KEYINPUT124), .B(G197gat), .Z(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n362_), .B(new_n413_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n846_), .A2(new_n680_), .A3(new_n901_), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n899_), .B(new_n900_), .S(new_n902_), .Z(G1352gat));
  AND2_X1   g702(.A1(new_n846_), .A2(new_n901_), .ZN(new_n904_));
  INV_X1    g703(.A(G204gat), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n904_), .B(new_n545_), .C1(KEYINPUT125), .C2(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n904_), .A2(new_n545_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT125), .B(G204gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1353gat));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910_));
  INV_X1    g709(.A(G211gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n585_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT126), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n804_), .A2(new_n405_), .A3(new_n901_), .A4(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n846_), .A2(new_n916_), .A3(new_n901_), .A4(new_n913_), .ZN(new_n917_));
  AND4_X1   g716(.A1(new_n910_), .A2(new_n915_), .A3(new_n911_), .A4(new_n917_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n915_), .A2(new_n917_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n904_), .A2(new_n921_), .A3(new_n593_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n904_), .A2(new_n634_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n921_), .ZN(G1355gat));
endmodule


