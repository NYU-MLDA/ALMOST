//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  AND4_X1   g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n206_), .A2(KEYINPUT80), .A3(new_n202_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n209_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n213_), .A2(new_n216_), .A3(new_n214_), .A4(new_n217_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(new_n223_), .A3(new_n219_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n226_), .A2(new_n227_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n227_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .A4(new_n209_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT4), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT89), .Z(new_n237_));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n225_), .A2(new_n228_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT92), .A4(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n229_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT91), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G57gat), .B(G85gat), .Z(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n248_), .B(KEYINPUT91), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n247_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n251_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n246_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n245_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n240_), .A2(new_n260_), .A3(new_n244_), .A4(new_n241_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT97), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(KEYINPUT97), .A3(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(G1gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT101), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G183gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT25), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .A4(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT78), .ZN(new_n281_));
  INV_X1    g080(.A(G169gat), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n284_), .A2(KEYINPUT24), .A3(new_n295_), .A4(new_n285_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n280_), .A2(new_n288_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n283_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n278_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n291_), .A2(new_n292_), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n295_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT79), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT30), .B(G99gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G43gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT31), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(G71gat), .Z(new_n311_));
  OR2_X1    g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G227gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n228_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n311_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n225_), .B2(KEYINPUT29), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n231_), .A2(new_n321_), .A3(new_n322_), .A4(new_n209_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G22gat), .B(G50gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n319_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n323_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT84), .A3(new_n325_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT21), .B1(new_n333_), .B2(KEYINPUT83), .ZN(new_n334_));
  INV_X1    g133(.A(G204gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G197gat), .ZN(new_n336_));
  INV_X1    g135(.A(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G204gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT83), .ZN(new_n339_));
  AND2_X1   g138(.A1(G211gat), .A2(G218gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n334_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n337_), .A2(G204gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n335_), .A2(G197gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT21), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n342_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n346_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AOI211_X1 g153(.A(KEYINPUT82), .B(new_n342_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n345_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n356_), .A2(KEYINPUT81), .B1(G228gat), .B2(G233gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT21), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT21), .B1(new_n336_), .B2(new_n338_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n353_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT82), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n352_), .A2(new_n346_), .A3(new_n353_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n344_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n357_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n356_), .A2(new_n358_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n328_), .A2(new_n332_), .A3(new_n367_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n331_), .A2(new_n325_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n357_), .A2(new_n366_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n370_), .A2(new_n371_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n319_), .B(new_n374_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n318_), .A2(new_n269_), .A3(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT18), .B(G64gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT98), .Z(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n297_), .A2(new_n304_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n365_), .A2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT87), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n399_));
  AOI21_X1  g198(.A(G176gat), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n303_), .A2(new_n295_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n274_), .A2(new_n279_), .A3(KEYINPUT85), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT85), .B1(new_n274_), .B2(new_n279_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n272_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n293_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n295_), .A2(KEYINPUT24), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n295_), .A2(KEYINPUT86), .A3(KEYINPUT24), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n284_), .A3(new_n285_), .A4(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT20), .B1(new_n356_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n394_), .B1(new_n414_), .B2(KEYINPUT95), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n400_), .A2(new_n401_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n411_), .A2(new_n294_), .A3(new_n288_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n405_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n419_), .B2(new_n365_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n392_), .B1(new_n415_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n419_), .B2(new_n365_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n416_), .B1(new_n365_), .B2(new_n393_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n356_), .A2(KEYINPUT88), .A3(new_n413_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(new_n391_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n389_), .B1(new_n423_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n394_), .A2(new_n391_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n428_), .A2(new_n391_), .B1(new_n431_), .B2(new_n420_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n388_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(KEYINPUT27), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(new_n391_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n420_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n437_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n433_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n436_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n384_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n388_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n229_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n261_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n434_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n263_), .A2(KEYINPUT93), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n263_), .B2(KEYINPUT93), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT94), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n439_), .A2(new_n440_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n451_), .A2(new_n452_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n448_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n433_), .A2(KEYINPUT32), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n423_), .B2(new_n429_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT96), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n432_), .A2(new_n459_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT96), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n464_), .B(new_n460_), .C1(new_n423_), .C2(new_n429_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n454_), .A2(new_n458_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n383_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT99), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n381_), .A2(new_n267_), .A3(new_n266_), .A4(new_n382_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n442_), .B2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n435_), .A2(new_n441_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n373_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n379_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n268_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(new_n475_), .A3(KEYINPUT99), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n318_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n443_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G29gat), .B(G36gat), .ZN(new_n483_));
  INV_X1    g282(.A(G50gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT72), .B(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  INV_X1    g290(.A(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n487_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n490_), .B1(new_n499_), .B2(new_n489_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT76), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n499_), .A2(new_n501_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n482_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n482_), .ZN(new_n507_));
  OAI221_X1 g306(.A(new_n507_), .B1(new_n501_), .B2(new_n499_), .C1(new_n500_), .C2(new_n503_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT100), .B1(new_n479_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT100), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n476_), .A2(new_n471_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n318_), .B1(new_n513_), .B2(new_n468_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n512_), .B(new_n509_), .C1(new_n514_), .C2(new_n443_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n520_), .A2(new_n521_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT67), .B(G71gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G78gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n523_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(KEYINPUT11), .A3(new_n522_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n535_));
  NAND2_X1  g334(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(KEYINPUT66), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT66), .B1(new_n535_), .B2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n534_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n543_), .A2(G99gat), .A3(G106gat), .A4(new_n537_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT7), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G85gat), .B(G92gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(KEYINPUT8), .A3(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(KEYINPUT8), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n534_), .B(KEYINPUT64), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT6), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT9), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G85gat), .A3(G92gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT10), .B(G99gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(G106gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n550_), .A2(new_n556_), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n559_), .A2(new_n560_), .B1(new_n547_), .B2(KEYINPUT8), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n553_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n533_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT69), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n563_), .B2(new_n533_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(KEYINPUT69), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n519_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI22_X1  g369(.A1(new_n533_), .A2(new_n563_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n533_), .A2(new_n563_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n533_), .B2(new_n563_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n572_), .B(new_n518_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT5), .B(G176gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G204gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n568_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n517_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n582_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n533_), .B(new_n497_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n592_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(new_n592_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n563_), .A2(new_n489_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n488_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT34), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n563_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT71), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n606_), .A2(new_n613_), .A3(new_n609_), .A4(new_n610_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n615_), .A2(KEYINPUT36), .A3(new_n616_), .A4(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n615_), .A2(KEYINPUT74), .A3(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n624_), .A3(new_n622_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT37), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n621_), .A2(new_n624_), .A3(new_n622_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n624_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n604_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n271_), .A2(new_n516_), .A3(new_n589_), .A4(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n588_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n271_), .B1(new_n635_), .B2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n270_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n585_), .A2(new_n587_), .A3(new_n509_), .A4(new_n603_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT102), .Z(new_n641_));
  NOR2_X1   g440(.A1(new_n630_), .A2(new_n631_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT103), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n479_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n641_), .A2(new_n645_), .A3(KEYINPUT104), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT104), .B1(new_n641_), .B2(new_n645_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n269_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT38), .B(new_n270_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n639_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n639_), .A2(new_n653_), .A3(new_n649_), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1324gat));
  NAND3_X1  g454(.A1(new_n641_), .A2(new_n645_), .A3(new_n442_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT106), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(G8gat), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(KEYINPUT106), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n493_), .B(new_n442_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n648_), .B2(new_n478_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT41), .Z(new_n667_));
  AND2_X1   g466(.A1(new_n635_), .A2(new_n633_), .ZN(new_n668_));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n318_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT108), .Z(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n383_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n668_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n648_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(new_n674_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n588_), .A2(new_n510_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n632_), .A2(new_n628_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n477_), .A2(new_n478_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n443_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n632_), .A2(new_n628_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n685_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n685_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n479_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n682_), .B(new_n604_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(KEYINPUT110), .A2(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n690_), .A3(new_n685_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n479_), .B2(new_n689_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n695_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n682_), .A3(new_n604_), .A4(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(new_n268_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G29gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n604_), .B1(new_n631_), .B2(new_n630_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT111), .Z(new_n705_));
  AOI211_X1 g504(.A(new_n588_), .B(new_n705_), .C1(new_n511_), .C2(new_n515_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n269_), .A2(G29gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n472_), .A2(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n706_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n705_), .ZN(new_n714_));
  AND4_X1   g513(.A1(new_n711_), .A2(new_n635_), .A3(new_n714_), .A4(new_n712_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n696_), .A2(new_n442_), .A3(new_n701_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n706_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n635_), .A2(new_n714_), .A3(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT112), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n721_), .A3(KEYINPUT45), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n718_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n716_), .A2(new_n718_), .A3(KEYINPUT46), .A4(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n696_), .A2(new_n318_), .A3(new_n701_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n478_), .A2(G43gat), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n728_), .A2(G43gat), .B1(new_n706_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g530(.A1(new_n696_), .A2(new_n674_), .A3(new_n701_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n674_), .A2(new_n484_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n732_), .A2(new_n484_), .B1(new_n707_), .B2(new_n734_), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n688_), .A2(new_n510_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n588_), .A3(new_n633_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n268_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n588_), .A2(new_n510_), .ZN(new_n741_));
  NOR4_X1   g540(.A1(new_n644_), .A2(new_n479_), .A3(new_n604_), .A4(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(G57gat), .A3(new_n268_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT115), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n740_), .A2(new_n744_), .ZN(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n442_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n442_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G64gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT48), .B(new_n746_), .C1(new_n742_), .C2(new_n442_), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n738_), .A2(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT116), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n742_), .B2(new_n318_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT49), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n318_), .A2(new_n754_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n738_), .B2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n742_), .B2(new_n674_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n739_), .A2(new_n759_), .A3(new_n674_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .ZN(G1335gat));
  AND2_X1   g567(.A1(new_n737_), .A2(new_n588_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n714_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n268_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n699_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n741_), .A2(new_n603_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n697_), .A2(KEYINPUT118), .A3(new_n698_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n269_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n771_), .B1(new_n777_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g577(.A(G92gat), .B1(new_n770_), .B2(new_n442_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n776_), .A2(new_n472_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n776_), .B2(new_n478_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n769_), .A2(new_n714_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n478_), .A2(new_n558_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT51), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n782_), .B(new_n787_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1338gat));
  OR2_X1    g588(.A1(new_n383_), .A2(G106gat), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n699_), .A2(new_n674_), .A3(new_n774_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G106gat), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n791_), .A3(G106gat), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n783_), .A2(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI221_X1 g596(.A(new_n797_), .B1(new_n793_), .B2(new_n794_), .C1(new_n783_), .C2(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  NAND2_X1  g598(.A1(new_n498_), .A2(new_n502_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n482_), .B(new_n800_), .C1(new_n500_), .C2(new_n502_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n508_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n574_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n575_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n571_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT55), .B1(new_n806_), .B2(new_n518_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n576_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n519_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n580_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n581_), .C1(new_n808_), .C2(new_n812_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n582_), .B(new_n803_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n810_), .B1(new_n809_), .B2(new_n519_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n576_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n580_), .B1(new_n822_), .B2(new_n811_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n815_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n583_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n803_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n819_), .A2(new_n828_), .A3(new_n690_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n509_), .A2(new_n582_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n802_), .B1(new_n586_), .B2(new_n582_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n642_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n642_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n829_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n589_), .A2(new_n633_), .A3(new_n510_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT54), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(KEYINPUT54), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n837_), .A2(new_n604_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n478_), .A2(new_n674_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n442_), .A2(new_n269_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n509_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n837_), .A2(new_n604_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n840_), .A2(new_n839_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n844_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT59), .B1(new_n853_), .B2(KEYINPUT121), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n852_), .B(new_n856_), .C1(KEYINPUT121), .C2(new_n853_), .ZN(new_n857_));
  AND4_X1   g656(.A1(new_n509_), .A2(new_n849_), .A3(new_n855_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n846_), .B1(new_n858_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n589_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n845_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  AND4_X1   g661(.A1(new_n588_), .A2(new_n849_), .A3(new_n855_), .A4(new_n857_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n854_), .B2(new_n604_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n867_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n604_), .A2(new_n865_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n849_), .A2(new_n855_), .A3(new_n857_), .A4(new_n870_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n869_), .A3(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n845_), .B2(new_n644_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT123), .B(G134gat), .ZN(new_n874_));
  AND4_X1   g673(.A1(new_n857_), .A2(new_n849_), .A3(new_n855_), .A4(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n690_), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n442_), .A2(new_n269_), .A3(new_n383_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n852_), .A2(new_n478_), .A3(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n510_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n589_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n212_), .ZN(G1345gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n604_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n878_), .A2(KEYINPUT124), .A3(new_n604_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n887_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n885_), .A3(new_n883_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(new_n878_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G162gat), .B1(new_n892_), .B2(new_n644_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n690_), .A2(G162gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT125), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(G1347gat));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n478_), .A2(new_n472_), .A3(new_n268_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(KEYINPUT126), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n674_), .B1(new_n898_), .B2(KEYINPUT126), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n852_), .A2(new_n509_), .A3(new_n900_), .A4(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(G169gat), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(G169gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n897_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n901_), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n841_), .A2(new_n510_), .A3(new_n899_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n397_), .A2(new_n399_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(new_n909_), .B2(new_n282_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(KEYINPUT62), .A3(new_n904_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n907_), .A2(new_n911_), .A3(new_n913_), .ZN(G1348gat));
  NOR3_X1   g713(.A1(new_n841_), .A2(new_n899_), .A3(new_n908_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n588_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G176gat), .ZN(G1349gat));
  AND2_X1   g716(.A1(new_n915_), .A2(new_n603_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n278_), .B2(new_n918_), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n272_), .A3(new_n644_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n915_), .A2(new_n690_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n301_), .ZN(G1351gat));
  NOR3_X1   g722(.A1(new_n841_), .A2(new_n318_), .A3(new_n472_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n475_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n510_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n337_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n589_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n335_), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n924_), .A2(new_n475_), .A3(new_n603_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n930_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n925_), .A2(new_n934_), .A3(new_n689_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n924_), .A2(new_n475_), .A3(new_n644_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(new_n936_), .ZN(G1355gat));
endmodule


