//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G85gat), .A3(G92gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G85gat), .B(G92gat), .ZN(new_n215_));
  OAI221_X1 g014(.A(new_n213_), .B1(new_n214_), .B2(G106gat), .C1(new_n212_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n215_), .B(KEYINPUT67), .Z(new_n221_));
  NOR2_X1   g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT7), .Z(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n210_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n221_), .B(new_n226_), .C1(new_n211_), .C2(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G43gat), .B(G50gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT15), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT75), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n218_), .A2(new_n219_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT35), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n236_), .A2(KEYINPUT73), .A3(new_n239_), .A4(new_n242_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(KEYINPUT35), .A3(new_n241_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(KEYINPUT35), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n244_), .B(new_n248_), .C1(new_n249_), .C2(KEYINPUT75), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n205_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT74), .B1(new_n247_), .B2(new_n250_), .ZN(new_n252_));
  OAI22_X1  g051(.A1(KEYINPUT36), .A2(new_n251_), .B1(new_n252_), .B2(new_n204_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT36), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n247_), .A2(new_n250_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n205_), .C1(new_n255_), .C2(KEYINPUT74), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT37), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G64gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G71gat), .B(G78gat), .ZN(new_n263_));
  OR3_X1    g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n263_), .A3(KEYINPUT11), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G15gat), .B(G22gat), .ZN(new_n267_));
  INV_X1    g066(.A(G1gat), .ZN(new_n268_));
  INV_X1    g067(.A(G8gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT14), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G1gat), .B(G8gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n266_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G127gat), .B(G155gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT16), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G183gat), .ZN(new_n280_));
  INV_X1    g079(.A(G211gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n277_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT76), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n277_), .A2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n287_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n258_), .A2(new_n259_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT96), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT0), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(G57gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(G57gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n296_), .A2(G85gat), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(G85gat), .B1(new_n296_), .B2(new_n297_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n304_), .A3(KEYINPUT1), .ZN(new_n305_));
  OR2_X1    g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n301_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n311_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n310_), .B(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n315_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n312_), .A2(new_n310_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n308_), .A2(new_n306_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n304_), .B1(new_n301_), .B2(KEYINPUT1), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n305_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n311_), .B(KEYINPUT3), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n310_), .B(KEYINPUT2), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n314_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n327_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n323_), .B(new_n324_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n313_), .A2(new_n341_), .A3(new_n320_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT91), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n321_), .A2(KEYINPUT91), .A3(new_n327_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n331_), .B1(new_n346_), .B2(KEYINPUT4), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n330_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n300_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT95), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n347_), .A2(new_n348_), .A3(new_n300_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT95), .B(new_n300_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT19), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT87), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT19), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n356_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n358_), .A2(new_n360_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT88), .ZN(new_n367_));
  INV_X1    g166(.A(new_n356_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n362_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G183gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT25), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT26), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G190gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n380_));
  AND3_X1   g179(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n379_), .A2(new_n380_), .A3(new_n383_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n382_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n371_), .A2(new_n375_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n384_), .A2(KEYINPUT22), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT22), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G169gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n396_), .A3(new_n385_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n397_), .A3(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT79), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n389_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  INV_X1    g202(.A(G204gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(G197gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(G197gat), .ZN(new_n406_));
  INV_X1    g205(.A(G197gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT21), .ZN(new_n410_));
  INV_X1    g209(.A(G218gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G211gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n281_), .A2(G218gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT85), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n405_), .A2(new_n408_), .A3(new_n410_), .A4(new_n406_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n404_), .A2(G197gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n407_), .A2(G204gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT21), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n400_), .A2(new_n402_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n426_));
  AND3_X1   g225(.A1(new_n409_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n417_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n387_), .B(KEYINPUT90), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n393_), .A2(new_n430_), .A3(new_n397_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n389_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n370_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n412_), .A2(new_n413_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n407_), .A2(G204gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n406_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(KEYINPUT21), .B2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n416_), .A2(new_n418_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n370_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT89), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n434_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G92gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G8gat), .B(G36gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT18), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n451_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n450_), .B(new_n451_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G64gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n455_), .A3(G92gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT32), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n448_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n442_), .A2(new_n443_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n389_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n401_), .B1(new_n389_), .B2(new_n398_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(new_n429_), .A3(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n431_), .A2(new_n389_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n439_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n466_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n439_), .A2(new_n470_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT20), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n467_), .A2(new_n468_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n473_), .B(new_n474_), .C1(new_n475_), .C2(new_n439_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n465_), .B1(KEYINPUT93), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n464_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n444_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n425_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n462_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n472_), .A2(new_n463_), .A3(new_n476_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n346_), .A2(new_n330_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n300_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n328_), .A2(new_n329_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n346_), .B2(KEYINPUT4), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n485_), .B(new_n486_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n492_));
  NOR4_X1   g291(.A1(new_n347_), .A2(new_n348_), .A3(new_n300_), .A4(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n353_), .A2(new_n492_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n355_), .A2(new_n481_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n336_), .A2(new_n339_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n429_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n429_), .A2(KEYINPUT83), .B1(G228gat), .B2(G233gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n498_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G22gat), .B(G50gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n504_), .A2(new_n505_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT86), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n504_), .A2(new_n505_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n503_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n506_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n509_), .A2(new_n515_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n502_), .B(new_n516_), .C1(new_n517_), .C2(new_n511_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n509_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n511_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n501_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n293_), .B1(new_n496_), .B2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT27), .B1(new_n485_), .B2(new_n486_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT27), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n458_), .A2(new_n526_), .A3(new_n461_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n448_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n486_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n472_), .A2(KEYINPUT99), .A3(new_n476_), .A4(new_n463_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT100), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n530_), .A2(new_n532_), .A3(KEYINPUT100), .A4(new_n533_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n524_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n355_), .A2(KEYINPUT97), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n352_), .B1(new_n350_), .B2(new_n349_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT97), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n354_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n538_), .A2(new_n539_), .A3(new_n542_), .A4(new_n522_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n518_), .A2(new_n521_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n540_), .A2(new_n354_), .B1(new_n480_), .B2(new_n478_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n492_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n352_), .A2(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n547_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n544_), .B(KEYINPUT96), .C1(new_n545_), .C2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n523_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n475_), .B(KEYINPUT30), .ZN(new_n551_));
  XOR2_X1   g350(.A(G71gat), .B(G99gat), .Z(new_n552_));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n551_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n555_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G15gat), .B(G43gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n341_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n558_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n550_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT101), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n550_), .A2(KEYINPUT101), .A3(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n539_), .A2(new_n542_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n544_), .A4(new_n538_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT64), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n238_), .A2(new_n266_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n573_), .B2(KEYINPUT68), .ZN(new_n574_));
  INV_X1    g373(.A(new_n266_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n229_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT68), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n573_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(KEYINPUT12), .A3(new_n573_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n238_), .A2(KEYINPUT12), .A3(new_n266_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n572_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT70), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(KEYINPUT71), .Z(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT13), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n235_), .A2(new_n273_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n273_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n232_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n273_), .B(new_n232_), .Z(new_n602_));
  INV_X1    g401(.A(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT77), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(G169gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n407_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT78), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n606_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n596_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n292_), .A2(new_n569_), .A3(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT102), .Z(new_n615_));
  INV_X1    g414(.A(new_n567_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n268_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n253_), .A2(new_n256_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n291_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n569_), .A2(new_n619_), .A3(new_n620_), .A4(new_n613_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT103), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n567_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n538_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n269_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G8gat), .B1(new_n621_), .B2(new_n538_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT39), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n623_), .B2(new_n561_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT104), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(KEYINPUT104), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(KEYINPUT41), .A3(new_n634_), .ZN(new_n638_));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n615_), .A2(new_n639_), .A3(new_n566_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(new_n638_), .A3(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n622_), .B2(new_n522_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n615_), .A2(new_n642_), .A3(new_n522_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n253_), .A2(new_n256_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n569_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n612_), .A2(new_n620_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n616_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(KEYINPUT37), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n569_), .A2(new_n653_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n569_), .A2(KEYINPUT105), .A3(new_n653_), .A4(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n569_), .A2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT43), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n649_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n652_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n663_), .C2(new_n649_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(G29gat), .A3(new_n616_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n651_), .B1(new_n669_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n650_), .A2(new_n673_), .A3(new_n626_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n626_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n649_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n653_), .B1(new_n569_), .B2(new_n656_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n658_), .B2(new_n657_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n679_), .B2(new_n660_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n680_), .B2(KEYINPUT44), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n664_), .A2(new_n652_), .A3(new_n665_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n675_), .B1(new_n683_), .B2(new_n673_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1329gat));
  AND2_X1   g485(.A1(new_n566_), .A2(G43gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n670_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G43gat), .B1(new_n650_), .B2(new_n566_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT107), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  INV_X1    g491(.A(new_n690_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(new_n693_), .C1(new_n668_), .C2(new_n688_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n691_), .A2(KEYINPUT47), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT47), .B1(new_n691_), .B2(new_n694_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n650_), .B2(new_n522_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n670_), .A2(G50gat), .A3(new_n522_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n669_), .B2(new_n699_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n596_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n292_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT108), .Z(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n611_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n569_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(G57gat), .A3(new_n567_), .ZN(new_n706_));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n569_), .A2(new_n619_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n596_), .A2(new_n611_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n708_), .A2(new_n291_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n710_), .B2(new_n616_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n706_), .A2(new_n711_), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n453_), .B1(new_n710_), .B2(new_n626_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n626_), .A2(new_n453_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n705_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT109), .Z(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n710_), .B2(new_n566_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NOR2_X1   g519(.A1(new_n561_), .A2(G71gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT110), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n705_), .B2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n710_), .B2(new_n522_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT50), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n522_), .A2(new_n724_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n705_), .B2(new_n727_), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n709_), .A2(new_n620_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n648_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G85gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n616_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n663_), .A2(new_n729_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n616_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n734_), .B2(new_n731_), .ZN(G1336gat));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n449_), .A3(new_n626_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n733_), .A2(new_n626_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n449_), .ZN(G1337gat));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n566_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n561_), .A2(new_n214_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n739_), .A2(G99gat), .B1(new_n730_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g541(.A(G106gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n663_), .A2(new_n522_), .A3(new_n729_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(KEYINPUT111), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n663_), .A2(new_n746_), .A3(new_n522_), .A4(new_n729_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n745_), .A2(KEYINPUT112), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT112), .B1(new_n745_), .B2(new_n747_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n730_), .A2(new_n743_), .A3(new_n522_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n744_), .A2(KEYINPUT111), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(G106gat), .A3(new_n747_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n756_), .B2(KEYINPUT52), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT53), .B1(new_n751_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n745_), .A2(KEYINPUT112), .A3(new_n747_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(KEYINPUT52), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n749_), .A2(new_n750_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n752_), .A4(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(G1339gat));
  NAND2_X1  g563(.A1(new_n611_), .A2(new_n589_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n579_), .A2(new_n572_), .A3(new_n580_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n581_), .B1(KEYINPUT55), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n572_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n590_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT56), .B(new_n590_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n605_), .A2(new_n609_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n599_), .A2(new_n603_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n597_), .A2(new_n777_), .B1(new_n602_), .B2(new_n600_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n609_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n592_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n619_), .B1(new_n774_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT115), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n772_), .A2(new_n773_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n765_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n647_), .B1(new_n787_), .B2(new_n780_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n784_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n589_), .A2(new_n779_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n654_), .A2(new_n655_), .B1(KEYINPUT58), .B2(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(KEYINPUT58), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n794_), .A2(new_n795_), .B1(new_n783_), .B2(new_n782_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n291_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n611_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n292_), .A2(KEYINPUT113), .A3(new_n799_), .A4(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n654_), .A2(new_n800_), .A3(new_n620_), .A4(new_n655_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT54), .B1(new_n802_), .B2(new_n803_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n798_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NOR4_X1   g608(.A1(new_n561_), .A2(new_n626_), .A3(new_n567_), .A4(new_n522_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(G113gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n611_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n793_), .A2(KEYINPUT58), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n656_), .A2(new_n795_), .A3(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n788_), .B2(KEYINPUT57), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n791_), .B1(new_n817_), .B2(KEYINPUT116), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n796_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n291_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n801_), .A2(new_n804_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n805_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n806_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n810_), .A2(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n811_), .A2(KEYINPUT59), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n611_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n814_), .B1(new_n830_), .B2(new_n813_), .ZN(G1340gat));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n812_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n832_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n829_), .A2(new_n701_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n812_), .A2(new_n837_), .A3(new_n620_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n829_), .A2(new_n620_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1342gat));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n829_), .B2(new_n656_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n811_), .A2(G134gat), .A3(new_n619_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n811_), .A2(KEYINPUT59), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(new_n828_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n656_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT117), .B(new_n846_), .C1(new_n849_), .C2(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n566_), .A2(new_n544_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n825_), .B2(new_n798_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n567_), .A2(new_n626_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n611_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n701_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n620_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(G162gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n856_), .A2(new_n864_), .A3(new_n647_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n854_), .A2(new_n656_), .A3(new_n855_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G162gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT118), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n870_), .A3(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n616_), .A2(new_n538_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n561_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n611_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT119), .Z(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n522_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n384_), .B1(new_n826_), .B2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n826_), .A2(new_n544_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n394_), .A2(new_n396_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n876_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1348gat));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n824_), .A2(new_n806_), .B1(new_n291_), .B2(new_n797_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n522_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n809_), .A2(KEYINPUT121), .A3(new_n544_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n874_), .A2(new_n596_), .A3(new_n385_), .A4(new_n561_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(KEYINPUT122), .A3(new_n890_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n826_), .A2(new_n544_), .A3(new_n701_), .A4(new_n875_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n385_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT120), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n898_), .A3(new_n385_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n893_), .A2(new_n894_), .B1(new_n897_), .B2(new_n899_), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n875_), .A2(new_n620_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n826_), .A2(new_n544_), .A3(new_n875_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n372_), .A2(new_n374_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n620_), .A2(new_n904_), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n902_), .A2(G183gat), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI221_X1 g707(.A(KEYINPUT123), .B1(new_n903_), .B2(new_n905_), .C1(new_n902_), .C2(G183gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1350gat));
  INV_X1    g709(.A(new_n656_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G190gat), .B1(new_n903_), .B2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n647_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n913_), .ZN(G1351gat));
  NAND3_X1  g713(.A1(new_n809_), .A2(new_n852_), .A3(new_n873_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT124), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n854_), .A2(new_n917_), .A3(new_n873_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n611_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g720(.A(new_n596_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n922_));
  AND2_X1   g721(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n924_), .ZN(G1353gat));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n917_), .B1(new_n854_), .B2(new_n873_), .ZN(new_n928_));
  NOR4_X1   g727(.A1(new_n886_), .A2(KEYINPUT124), .A3(new_n853_), .A4(new_n874_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n620_), .B(new_n927_), .C1(new_n928_), .C2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT126), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n919_), .A2(new_n932_), .A3(new_n620_), .A4(new_n927_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n620_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n931_), .A2(new_n933_), .A3(new_n936_), .ZN(G1354gat));
  AOI21_X1  g736(.A(G218gat), .B1(new_n919_), .B2(new_n647_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n656_), .A2(G218gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT127), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n919_), .B2(new_n940_), .ZN(G1355gat));
endmodule


