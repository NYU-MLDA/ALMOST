//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT13), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(KEYINPUT13), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(KEYINPUT9), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(KEYINPUT9), .B2(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n215_), .B2(new_n216_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n212_), .B(new_n214_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT8), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(KEYINPUT8), .ZN(new_n224_));
  OAI22_X1  g023(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  OR4_X1    g024(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n214_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n209_), .A2(new_n210_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n206_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT68), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n231_), .A3(new_n206_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n223_), .B(new_n224_), .C1(new_n227_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n214_), .A2(new_n226_), .A3(new_n225_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n222_), .A3(KEYINPUT8), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n234_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n221_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n244_));
  XOR2_X1   g043(.A(G71gat), .B(G78gat), .Z(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT12), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G230gat), .A2(G233gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n221_), .A2(new_n234_), .A3(new_n237_), .A4(new_n248_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT12), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n234_), .A2(new_n237_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n221_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n249_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n254_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n253_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT70), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n265_), .A3(new_n262_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT73), .B(G120gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n270_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n260_), .A2(new_n264_), .A3(new_n266_), .A4(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n204_), .B(new_n205_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n276_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT13), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(KEYINPUT75), .A3(new_n278_), .A4(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G15gat), .B(G22gat), .Z(new_n288_));
  NAND2_X1  g087(.A1(G1gat), .A2(G8gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(KEYINPUT14), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT79), .ZN(new_n291_));
  XOR2_X1   g090(.A(G1gat), .B(G8gat), .Z(new_n292_));
  AND2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G229gat), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n299_), .B(KEYINPUT15), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n295_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G141gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G169gat), .B(G197gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n305_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n287_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT89), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n318_), .B(new_n319_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT89), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT31), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT88), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G71gat), .B(G99gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(KEYINPUT85), .A2(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(KEYINPUT85), .A2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330_));
  INV_X1    g129(.A(G169gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n328_), .A2(new_n329_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT83), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT86), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(KEYINPUT23), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n343_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n345_), .B1(KEYINPUT86), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  INV_X1    g149(.A(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n337_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n350_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT25), .B1(new_n350_), .B2(KEYINPUT82), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n336_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n339_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n344_), .A2(new_n338_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT24), .ZN(new_n365_));
  INV_X1    g164(.A(G176gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n331_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n361_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n369_));
  AOI211_X1 g168(.A(KEYINPUT84), .B(new_n369_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n358_), .B(new_n360_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n354_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n326_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G15gat), .B(G43gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n375_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT18), .B(G64gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT19), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n367_), .B1(new_n336_), .B2(new_n359_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n356_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n340_), .A2(KEYINPUT23), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n338_), .A2(KEYINPUT83), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n344_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n394_), .B2(new_n346_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n390_), .B1(new_n395_), .B2(new_n345_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n335_), .A2(KEYINPUT96), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT96), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT97), .B1(new_n334_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n364_), .A2(new_n352_), .ZN(new_n402_));
  AND2_X1   g201(.A1(KEYINPUT85), .A2(G176gat), .ZN(new_n403_));
  AND2_X1   g202(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n327_), .A2(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n401_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G197gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(G204gat), .ZN(new_n411_));
  INV_X1    g210(.A(G204gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(G197gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT21), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(G197gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(G204gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT21), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n419_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n416_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT21), .A3(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n396_), .A2(new_n409_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT20), .ZN(new_n426_));
  INV_X1    g225(.A(new_n424_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n426_), .A2(KEYINPUT100), .B1(new_n372_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n429_), .A3(KEYINPUT20), .ZN(new_n430_));
  AOI211_X1 g229(.A(KEYINPUT101), .B(new_n387_), .C1(new_n428_), .C2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT101), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(KEYINPUT100), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n372_), .A2(new_n427_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n430_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n435_), .B2(new_n386_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n354_), .A2(new_n371_), .A3(new_n424_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n409_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n401_), .A2(new_n402_), .A3(new_n408_), .A4(KEYINPUT98), .ZN(new_n441_));
  INV_X1    g240(.A(new_n349_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n440_), .A2(new_n441_), .B1(new_n442_), .B2(new_n390_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT20), .B(new_n438_), .C1(new_n443_), .C2(new_n424_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(new_n386_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n384_), .B1(new_n437_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n386_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n441_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n424_), .A3(new_n396_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n434_), .A3(KEYINPUT20), .A4(new_n387_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n450_), .A3(new_n384_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT27), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT103), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT27), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n447_), .A2(new_n450_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(new_n384_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n451_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n435_), .A2(new_n386_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT101), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n435_), .A2(new_n432_), .A3(new_n386_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n445_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n384_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT103), .ZN(new_n466_));
  INV_X1    g265(.A(new_n452_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n453_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G141gat), .ZN(new_n470_));
  INV_X1    g269(.A(G148gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT90), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT3), .ZN(new_n473_));
  NAND3_X1  g272(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(new_n470_), .A3(new_n471_), .A4(KEYINPUT90), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT2), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .A4(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n470_), .A2(new_n471_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n480_), .A2(KEYINPUT1), .B1(new_n470_), .B2(new_n471_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n322_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT4), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n479_), .A2(new_n482_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n321_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(KEYINPUT4), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT99), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n490_), .A2(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n495_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n491_), .A2(new_n494_), .A3(KEYINPUT99), .A4(new_n496_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n209_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT0), .B(G57gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G78gat), .B(G106gat), .Z(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n514_));
  INV_X1    g313(.A(G228gat), .ZN(new_n515_));
  INV_X1    g314(.A(G233gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n514_), .A2(new_n424_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n489_), .A2(KEYINPUT92), .A3(KEYINPUT29), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n492_), .B2(new_n513_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n522_), .A3(new_n427_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n523_), .A2(KEYINPUT93), .A3(new_n517_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT93), .B1(new_n523_), .B2(new_n517_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n512_), .B(new_n519_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n492_), .A2(new_n513_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G22gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n527_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n427_), .B1(new_n514_), .B2(KEYINPUT92), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n492_), .A2(new_n521_), .A3(new_n513_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n517_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n523_), .A2(KEYINPUT93), .A3(new_n517_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n518_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(new_n512_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n532_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n539_), .B2(new_n512_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n512_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT95), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n526_), .A2(KEYINPUT94), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n537_), .A2(new_n538_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n512_), .A4(new_n519_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n543_), .A2(new_n546_), .A3(new_n547_), .A4(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n531_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n541_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n469_), .A2(new_n511_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n463_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT102), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n456_), .A2(new_n556_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT102), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n463_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n559_), .A2(new_n511_), .A3(new_n560_), .A4(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n457_), .A2(new_n458_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n510_), .B(KEYINPUT33), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n491_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n500_), .A2(new_n496_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n507_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n555_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n380_), .B1(new_n554_), .B2(new_n570_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT103), .B(new_n452_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n466_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(KEYINPUT104), .A3(new_n553_), .A4(new_n459_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n453_), .A2(new_n553_), .A3(new_n459_), .A4(new_n468_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT104), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n511_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n575_), .A2(new_n578_), .A3(new_n579_), .A4(new_n379_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n317_), .B1(new_n571_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n241_), .A2(new_n306_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n221_), .A2(new_n234_), .A3(new_n237_), .A4(new_n299_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT76), .B(KEYINPUT35), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n586_), .B(new_n588_), .C1(new_n583_), .C2(KEYINPUT77), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n582_), .A2(new_n591_), .A3(new_n583_), .A4(new_n589_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n593_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n593_), .A2(new_n599_), .B1(new_n597_), .B2(new_n596_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT78), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n593_), .A2(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n596_), .A2(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n593_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(KEYINPUT78), .A3(KEYINPUT37), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT81), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT17), .Z(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n248_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n295_), .B(new_n620_), .Z(new_n621_));
  OR2_X1    g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(KEYINPUT17), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n611_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n581_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(G1gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n511_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT38), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(new_n609_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n581_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(new_n511_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n629_), .B2(new_n634_), .ZN(G1324gat));
  INV_X1    g434(.A(G8gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n636_), .A3(new_n469_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n469_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(G8gat), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n638_), .B2(G8gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n628_), .A2(new_n645_), .A3(new_n379_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n633_), .B2(new_n379_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n633_), .B2(new_n555_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n628_), .A2(new_n652_), .A3(new_n555_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(new_n609_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n625_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n581_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n511_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n604_), .A2(new_n610_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n571_), .B2(new_n580_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n317_), .A2(new_n625_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT44), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G29gat), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n579_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n571_), .A2(new_n580_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n664_), .B1(new_n670_), .B2(new_n611_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT43), .B(new_n662_), .C1(new_n571_), .C2(new_n580_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT44), .B(new_n666_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n661_), .B1(new_n669_), .B2(new_n673_), .ZN(G1328gat));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n469_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G36gat), .B1(new_n667_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n469_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n659_), .A2(G36gat), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT46), .B1(new_n681_), .B2(KEYINPUT108), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n683_), .B(new_n684_), .C1(new_n676_), .C2(new_n680_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1329gat));
  NAND3_X1  g485(.A1(new_n673_), .A2(G43gat), .A3(new_n379_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n659_), .A2(new_n380_), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n687_), .A2(new_n667_), .B1(G43gat), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g489(.A1(new_n673_), .A2(G50gat), .A3(new_n555_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n659_), .A2(new_n553_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n691_), .A2(new_n667_), .B1(G50gat), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT109), .ZN(G1331gat));
  AOI21_X1  g493(.A(new_n316_), .B1(new_n571_), .B2(new_n580_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n287_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n632_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n579_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n695_), .B(KEYINPUT111), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(new_n627_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n511_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n699_), .B1(new_n707_), .B2(new_n698_), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n697_), .B2(new_n677_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(new_n706_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n677_), .A2(G64gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(G1333gat));
  OAI21_X1  g512(.A(G71gat), .B1(new_n697_), .B2(new_n380_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n380_), .A2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n711_), .B2(new_n716_), .ZN(G1334gat));
  OAI21_X1  g516(.A(G78gat), .B1(new_n697_), .B2(new_n553_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT50), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n553_), .A2(G78gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n711_), .B2(new_n720_), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n287_), .A2(new_n316_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n626_), .B(new_n722_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(new_n209_), .A3(new_n579_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n700_), .A2(new_n696_), .A3(new_n658_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(new_n579_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(new_n209_), .ZN(G1336gat));
  NOR3_X1   g526(.A1(new_n723_), .A2(new_n210_), .A3(new_n677_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n725_), .A2(new_n677_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n210_), .ZN(G1337gat));
  OAI21_X1  g529(.A(G99gat), .B1(new_n723_), .B2(new_n380_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n379_), .A2(new_n215_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n725_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n665_), .A2(new_n555_), .A3(new_n626_), .A4(new_n722_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n735_), .B(G106gat), .C1(new_n723_), .C2(new_n553_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n555_), .A2(new_n216_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n737_), .A2(new_n739_), .B1(new_n725_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  OAI221_X1 g542(.A(new_n743_), .B1(new_n725_), .B2(new_n740_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  NAND2_X1  g544(.A1(new_n662_), .A2(new_n625_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n316_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n281_), .A2(new_n747_), .A3(new_n286_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT54), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n287_), .A2(new_n627_), .A3(new_n750_), .A4(new_n747_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n253_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n260_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n252_), .A2(KEYINPUT55), .A3(new_n253_), .A4(new_n259_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n758_), .B2(new_n274_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT56), .B(new_n273_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n277_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n279_), .A2(new_n280_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n302_), .A2(new_n303_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n300_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n312_), .A3(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n315_), .A2(new_n766_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n762_), .A2(new_n316_), .B1(new_n763_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n609_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n768_), .B2(new_n609_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n758_), .A2(new_n274_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT56), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n758_), .A2(new_n753_), .A3(new_n274_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(new_n277_), .A3(new_n767_), .A4(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n777_), .B1(new_n610_), .B2(new_n604_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT114), .B1(new_n776_), .B2(new_n777_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n762_), .A2(new_n780_), .A3(KEYINPUT58), .A4(new_n767_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n772_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n752_), .B1(new_n783_), .B2(new_n626_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n575_), .A2(new_n578_), .A3(new_n511_), .A4(new_n379_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n316_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n784_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(KEYINPUT115), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n785_), .A2(KEYINPUT115), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n768_), .A2(new_n769_), .A3(new_n609_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n772_), .A2(new_n782_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n772_), .A2(new_n782_), .A3(KEYINPUT116), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n625_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n790_), .B(new_n791_), .C1(new_n797_), .C2(new_n752_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n789_), .B1(new_n798_), .B2(new_n788_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n747_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n787_), .B1(new_n800_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n287_), .B2(G120gat), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n786_), .B(new_n803_), .C1(new_n802_), .C2(G120gat), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G120gat), .B1(new_n799_), .B2(new_n287_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1341gat));
  AOI21_X1  g607(.A(KEYINPUT118), .B1(new_n625_), .B2(G127gat), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n625_), .B(new_n786_), .C1(new_n799_), .C2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n799_), .A2(KEYINPUT118), .A3(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(G1342gat));
  XNOR2_X1  g612(.A(KEYINPUT119), .B(G134gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n799_), .A2(new_n662_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G134gat), .B1(new_n786_), .B2(new_n609_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1343gat));
  NOR2_X1   g616(.A1(new_n784_), .A2(new_n379_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(new_n511_), .A3(new_n555_), .A4(new_n677_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n747_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(new_n470_), .ZN(G1344gat));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n287_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT120), .B(G148gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  NOR2_X1   g623(.A1(new_n819_), .A2(new_n626_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT61), .B(G155gat), .Z(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  NAND2_X1  g626(.A1(new_n611_), .A2(G162gat), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT122), .Z(new_n829_));
  NOR2_X1   g628(.A1(new_n819_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n819_), .B2(new_n657_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT121), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n831_), .C1(new_n819_), .C2(new_n657_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n830_), .B1(new_n833_), .B2(new_n835_), .ZN(G1347gat));
  NAND2_X1  g635(.A1(new_n749_), .A2(new_n751_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n793_), .A2(new_n794_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n838_), .A2(new_n770_), .A3(new_n796_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n839_), .B2(new_n625_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n677_), .A2(new_n511_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n379_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n555_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n840_), .A2(new_n841_), .A3(new_n316_), .A4(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n316_), .B(new_n844_), .C1(new_n797_), .C2(new_n752_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n847_), .A3(G169gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n797_), .A2(new_n752_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n844_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n316_), .C1(new_n405_), .C2(new_n404_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n845_), .A2(new_n847_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n854_), .A3(new_n855_), .ZN(G1348gat));
  OAI21_X1  g655(.A(KEYINPUT124), .B1(new_n784_), .B2(new_n555_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n626_), .B1(new_n793_), .B2(new_n792_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n837_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n553_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n843_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n287_), .A2(new_n366_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n857_), .A2(new_n861_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n851_), .A2(new_n287_), .A3(new_n852_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n328_), .A2(new_n329_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT125), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n864_), .B(new_n870_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1349gat));
  NAND4_X1  g671(.A1(new_n857_), .A2(new_n861_), .A3(new_n625_), .A4(new_n862_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n626_), .A2(new_n389_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n873_), .A2(new_n350_), .B1(new_n853_), .B2(new_n874_), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n853_), .A2(new_n356_), .A3(new_n609_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n851_), .A2(new_n662_), .A3(new_n852_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n351_), .B2(new_n877_), .ZN(G1351gat));
  NOR3_X1   g677(.A1(new_n677_), .A2(new_n511_), .A3(new_n553_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n818_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n747_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n410_), .ZN(G1352gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n287_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT126), .B(G204gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1353gat));
  NOR2_X1   g684(.A1(new_n880_), .A2(new_n626_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n886_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT63), .B(G211gat), .Z(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(new_n888_), .ZN(G1354gat));
  INV_X1    g688(.A(new_n880_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n890_), .A2(G218gat), .A3(new_n611_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G218gat), .B1(new_n890_), .B2(new_n609_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1355gat));
endmodule


