//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  NAND2_X1  g000(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(KEYINPUT75), .A3(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G183gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT76), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n205_), .A4(new_n203_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT77), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT24), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n230_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n216_), .A2(new_n229_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G169gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT81), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(KEYINPUT81), .A3(G169gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n218_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT22), .B1(KEYINPUT80), .B2(G169gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT82), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  AOI21_X1  g049(.A(G176gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .A4(new_n244_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n225_), .A2(new_n227_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n237_), .A2(new_n231_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n239_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G15gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n260_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT31), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G43gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G134gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G127gat), .ZN(new_n270_));
  INV_X1    g069(.A(G127gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G134gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G120gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G113gat), .ZN(new_n275_));
  INV_X1    g074(.A(G113gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G120gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n270_), .A2(new_n272_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n268_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n264_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G233gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT87), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(KEYINPUT87), .ZN(new_n287_));
  OAI21_X1  g086(.A(G228gat), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G197gat), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G197gat), .A2(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(KEYINPUT21), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  INV_X1    g104(.A(G141gat), .ZN(new_n306_));
  INV_X1    g105(.A(G148gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT84), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n315_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n309_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n315_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n325_), .B(new_n326_), .C1(new_n327_), .C2(KEYINPUT1), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n304_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n289_), .B1(new_n303_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n322_), .A2(new_n328_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT88), .B1(new_n299_), .B2(new_n300_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n288_), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT89), .Z(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n340_));
  XOR2_X1   g139(.A(G22gat), .B(G50gat), .Z(new_n341_));
  NAND4_X1  g140(.A1(new_n322_), .A2(new_n328_), .A3(new_n304_), .A4(new_n338_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n335_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n336_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n337_), .B1(new_n351_), .B2(KEYINPUT90), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n330_), .A2(new_n334_), .A3(new_n353_), .A4(new_n336_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n343_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n341_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT86), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n346_), .A2(new_n359_), .A3(new_n343_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n350_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n237_), .B2(new_n231_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT26), .B(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n213_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT24), .A4(new_n224_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n256_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n241_), .A2(new_n370_), .A3(new_n218_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n228_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n368_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT20), .B1(new_n373_), .B2(new_n301_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n299_), .A2(new_n300_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n239_), .B2(new_n259_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT19), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n374_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n378_), .B(KEYINPUT91), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n373_), .B2(new_n301_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n239_), .A2(new_n259_), .A3(new_n375_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n380_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT97), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n388_), .A2(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n389_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(KEYINPUT97), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n379_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n384_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n391_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n390_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n374_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n260_), .A2(new_n301_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n378_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n384_), .A2(new_n385_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n381_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n390_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT27), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n362_), .A2(new_n402_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n331_), .A2(new_n282_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(KEYINPUT4), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n322_), .A2(new_n281_), .A3(new_n328_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n281_), .B1(new_n328_), .B2(new_n322_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n421_), .B2(KEYINPUT4), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n322_), .A2(new_n281_), .A3(new_n328_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n415_), .A2(new_n418_), .A3(KEYINPUT4), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n417_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G85gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT0), .B(G57gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n419_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(KEYINPUT94), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n415_), .A2(KEYINPUT4), .A3(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT92), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n416_), .B1(new_n437_), .B2(new_n424_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n430_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n435_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n431_), .B1(new_n438_), .B2(new_n432_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT95), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n431_), .C1(new_n438_), .C2(new_n432_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT96), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT96), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n442_), .A2(new_n444_), .A3(new_n449_), .A4(new_n446_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n412_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n362_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n380_), .A2(new_n453_), .A3(new_n386_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n398_), .A2(new_n399_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n447_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n409_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(new_n391_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n414_), .B1(new_n420_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT93), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT93), .B(new_n461_), .C1(new_n422_), .C2(new_n425_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n430_), .B1(new_n421_), .B2(new_n414_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n426_), .A2(KEYINPUT33), .A3(new_n433_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n459_), .A2(new_n467_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n452_), .B1(new_n457_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n284_), .B1(new_n451_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n448_), .A2(new_n450_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(new_n284_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n402_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n411_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n362_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT98), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n402_), .A2(new_n411_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT98), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n362_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n473_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G183gat), .B(G211gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n487_), .A2(KEYINPUT11), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT70), .ZN(new_n497_));
  INV_X1    g296(.A(G15gat), .ZN(new_n498_));
  INV_X1    g297(.A(G22gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G15gat), .A2(G22gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G1gat), .A2(G8gat), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n500_), .A2(new_n501_), .B1(KEYINPUT14), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n497_), .B(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n495_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n495_), .A2(new_n504_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G127gat), .B(G155gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n511_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n486_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n486_), .A3(new_n513_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n517_), .A3(new_n507_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n516_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n514_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n521_), .B2(KEYINPUT17), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT67), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT15), .Z(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT10), .B(G99gat), .Z(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G85gat), .B(G92gat), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT9), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT6), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(G85gat), .A3(G92gat), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n534_), .A2(new_n536_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT7), .ZN(new_n546_));
  INV_X1    g345(.A(G99gat), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n533_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n545_), .B(new_n548_), .C1(new_n538_), .C2(new_n540_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n535_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n549_), .B2(new_n535_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n531_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n527_), .B1(new_n555_), .B2(KEYINPUT68), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n530_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n560_), .A3(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT36), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n563_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(KEYINPUT100), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(KEYINPUT100), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n485_), .A2(new_n522_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n492_), .A2(new_n491_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n488_), .A2(new_n489_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n553_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n493_), .B(new_n544_), .C1(new_n552_), .C2(new_n551_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT64), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT65), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT12), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n553_), .A2(new_n591_), .A3(new_n581_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n589_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT65), .B(new_n587_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n588_), .B(new_n602_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(KEYINPUT66), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT66), .B1(new_n601_), .B2(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n578_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(KEYINPUT13), .A3(new_n604_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G113gat), .B(G141gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT74), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n504_), .B(new_n530_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(KEYINPUT73), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT73), .B1(new_n615_), .B2(new_n617_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n531_), .A2(new_n504_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n504_), .A2(new_n530_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n617_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n614_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n614_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n626_), .B(new_n627_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT99), .B1(new_n610_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n632_));
  INV_X1    g431(.A(new_n629_), .ZN(new_n633_));
  AOI211_X1 g432(.A(new_n632_), .B(new_n633_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n577_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(KEYINPUT101), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n630_), .A2(new_n634_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n577_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n474_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n457_), .A2(new_n471_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n362_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n412_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n647_), .A2(new_n284_), .B1(new_n483_), .B2(new_n475_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n633_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT69), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT37), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT37), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n572_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n569_), .A2(new_n650_), .A3(KEYINPUT37), .A4(new_n571_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n610_), .A2(new_n522_), .A3(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(G1gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n474_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT38), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n643_), .A2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(G8gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n480_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n658_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n636_), .A2(KEYINPUT102), .A3(new_n480_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n663_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n636_), .B2(new_n480_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT40), .B(new_n665_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  INV_X1    g475(.A(new_n284_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n658_), .A2(new_n498_), .A3(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n679_), .B2(G15gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1326gat));
  NAND3_X1  g481(.A1(new_n658_), .A2(new_n499_), .A3(new_n452_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n452_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G22gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G22gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT103), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1327gat));
  OR2_X1    g491(.A1(new_n522_), .A2(new_n572_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n610_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n649_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n474_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n630_), .A2(new_n634_), .A3(new_n522_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n656_), .B1(new_n485_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n648_), .A2(KEYINPUT104), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n655_), .A2(new_n699_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT105), .B1(new_n648_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n485_), .A2(new_n706_), .A3(new_n699_), .A4(new_n655_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n698_), .B1(new_n703_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n698_), .B(KEYINPUT44), .C1(new_n703_), .C2(new_n708_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n474_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n697_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n664_), .A3(new_n712_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n480_), .B(KEYINPUT106), .Z(new_n720_));
  NAND4_X1  g519(.A1(new_n695_), .A2(new_n649_), .A3(new_n719_), .A4(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT45), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n716_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n722_), .B1(new_n717_), .B2(G36gat), .ZN(new_n727_));
  INV_X1    g526(.A(new_n716_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(KEYINPUT107), .A3(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1329gat));
  NAND4_X1  g529(.A1(new_n711_), .A2(G43gat), .A3(new_n677_), .A4(new_n712_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n696_), .A2(new_n677_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(G43gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n696_), .B2(new_n452_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n452_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n713_), .B2(new_n737_), .ZN(G1331gat));
  NAND3_X1  g537(.A1(new_n577_), .A2(new_n633_), .A3(new_n694_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n642_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n485_), .B2(new_n633_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n610_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n485_), .A2(KEYINPUT110), .A3(new_n633_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n522_), .A3(new_n656_), .A4(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n642_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n748_), .B2(new_n747_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n741_), .B1(new_n750_), .B2(new_n740_), .ZN(G1332gat));
  INV_X1    g550(.A(G64gat), .ZN(new_n752_));
  INV_X1    g551(.A(new_n739_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n720_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT48), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n720_), .A2(new_n752_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT113), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n747_), .B2(new_n757_), .ZN(G1333gat));
  OAI21_X1  g557(.A(G71gat), .B1(new_n739_), .B2(new_n284_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT49), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n284_), .A2(G71gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n747_), .B2(new_n761_), .ZN(G1334gat));
  OAI21_X1  g561(.A(G78gat), .B1(new_n739_), .B2(new_n362_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT50), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n362_), .A2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n747_), .B2(new_n765_), .ZN(G1335gat));
  OR2_X1    g565(.A1(new_n703_), .A2(new_n708_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n522_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n694_), .A2(new_n633_), .A3(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT114), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n474_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G85gat), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n743_), .A2(new_n744_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n693_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n642_), .A2(G85gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1336gat));
  INV_X1    g577(.A(new_n776_), .ZN(new_n779_));
  INV_X1    g578(.A(G92gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n664_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n771_), .A2(new_n720_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n780_), .ZN(G1337gat));
  AND3_X1   g582(.A1(new_n779_), .A2(new_n532_), .A3(new_n677_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n547_), .B1(new_n771_), .B2(new_n677_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n784_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n533_), .A3(new_n452_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n767_), .A2(new_n452_), .A3(new_n770_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n791_), .B(new_n798_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  AOI21_X1  g599(.A(new_n627_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n623_), .A2(new_n616_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n622_), .B2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n603_), .A2(new_n628_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n593_), .A2(new_n586_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT65), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n593_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n587_), .A2(KEYINPUT116), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n593_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n593_), .A2(new_n809_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n587_), .A2(KEYINPUT55), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n600_), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n815_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT58), .B(new_n804_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n655_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n814_), .A2(new_n815_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n815_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT58), .B1(new_n822_), .B2(new_n804_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n629_), .B(new_n603_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n608_), .A2(new_n628_), .A3(new_n604_), .A4(new_n803_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n825_), .A2(new_n826_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n629_), .A2(new_n603_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n628_), .A2(new_n803_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n605_), .A2(new_n606_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n572_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n828_), .A3(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n610_), .A2(new_n656_), .A3(new_n633_), .A4(new_n522_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n836_), .A2(new_n768_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n483_), .A2(new_n474_), .A3(new_n677_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT117), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n629_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n842_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n838_), .A2(new_n839_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n827_), .A2(KEYINPUT57), .B1(new_n819_), .B2(new_n823_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n833_), .A2(new_n834_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n768_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT118), .B(new_n768_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n847_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n845_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n276_), .B1(new_n629_), .B2(KEYINPUT119), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(KEYINPUT119), .B2(new_n276_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n844_), .B1(new_n857_), .B2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(new_n274_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n843_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n274_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT120), .ZN(new_n863_));
  OAI21_X1  g662(.A(G120gat), .B1(new_n856_), .B2(new_n610_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n856_), .B2(new_n768_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n843_), .A2(new_n271_), .A3(new_n522_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1342gat));
  NOR2_X1   g667(.A1(new_n656_), .A2(new_n269_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n845_), .B(new_n869_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n840_), .A2(new_n576_), .A3(new_n842_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT121), .B1(new_n871_), .B2(G134gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n850_), .A2(new_n846_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n842_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n873_), .B(new_n269_), .C1(new_n876_), .C2(new_n576_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n870_), .A2(new_n872_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n870_), .A2(new_n872_), .A3(KEYINPUT122), .A4(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n677_), .A2(new_n362_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n874_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n720_), .A2(new_n642_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n633_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n306_), .ZN(G1344gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n610_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT123), .B(G148gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1345gat));
  NAND4_X1  g690(.A1(new_n874_), .A2(new_n522_), .A3(new_n883_), .A4(new_n885_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT124), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(KEYINPUT124), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n886_), .B2(new_n656_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n576_), .A2(G162gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n886_), .B2(new_n900_), .ZN(G1347gat));
  INV_X1    g700(.A(new_n853_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT118), .B1(new_n836_), .B2(new_n768_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n846_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n720_), .A2(new_n642_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n284_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n904_), .A2(new_n629_), .A3(new_n362_), .A4(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G169gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n907_), .A2(G169gat), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n241_), .A2(new_n370_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n907_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n910_), .A2(new_n912_), .A3(new_n914_), .ZN(G1348gat));
  NOR2_X1   g714(.A1(new_n854_), .A2(new_n452_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n694_), .A3(new_n906_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n840_), .A2(new_n452_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n906_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n919_), .A2(new_n218_), .A3(new_n610_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n917_), .A2(new_n218_), .B1(new_n918_), .B2(new_n920_), .ZN(G1349gat));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n768_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G183gat), .B1(new_n918_), .B2(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n919_), .A2(new_n768_), .A3(new_n213_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n916_), .B2(new_n924_), .ZN(G1350gat));
  NAND2_X1  g724(.A1(new_n916_), .A2(new_n906_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G190gat), .B1(new_n926_), .B2(new_n656_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n575_), .A2(new_n365_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1351gat));
  INV_X1    g728(.A(new_n905_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n884_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n633_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n293_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n610_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n294_), .ZN(G1353gat));
  AOI21_X1  g734(.A(new_n768_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n874_), .A2(new_n883_), .A3(new_n930_), .A4(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n938_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n939_), .B2(new_n941_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n931_), .B2(new_n656_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n576_), .A2(G218gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n931_), .B2(new_n946_), .ZN(G1355gat));
endmodule


