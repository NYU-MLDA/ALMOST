//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT64), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT64), .B1(new_n203_), .B2(new_n205_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(KEYINPUT9), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n208_), .B(new_n213_), .C1(G106gat), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n203_), .A2(new_n205_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n217_), .A2(new_n218_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n212_), .ZN(new_n226_));
  OAI211_X1 g025(.A(KEYINPUT67), .B(KEYINPUT8), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n206_), .A2(new_n207_), .A3(new_n224_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n207_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n224_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT64), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n236_), .A2(KEYINPUT65), .A3(new_n230_), .A4(new_n212_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n218_), .A2(new_n224_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n203_), .A2(new_n205_), .A3(new_n216_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n212_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n242_), .B2(KEYINPUT8), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n215_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G78gat), .ZN(new_n248_));
  INV_X1    g047(.A(G78gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n249_), .A3(new_n246_), .ZN(new_n250_));
  INV_X1    g049(.A(G64gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G57gat), .ZN(new_n252_));
  INV_X1    g051(.A(G57gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G64gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT11), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT11), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(new_n250_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n250_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n249_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n255_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n244_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n215_), .B(new_n266_), .C1(new_n238_), .C2(new_n243_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G230gat), .A2(G233gat), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(KEYINPUT12), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT73), .B1(new_n244_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n226_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n230_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n227_), .A3(new_n232_), .A4(new_n237_), .ZN(new_n281_));
  AOI211_X1 g080(.A(new_n277_), .B(new_n274_), .C1(new_n281_), .C2(new_n215_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n270_), .B(new_n273_), .C1(new_n276_), .C2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(KEYINPUT71), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n244_), .A2(new_n286_), .A3(new_n267_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n271_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n281_), .A2(KEYINPUT70), .A3(new_n215_), .A4(new_n266_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n285_), .A2(new_n287_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n272_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(KEYINPUT72), .A3(new_n292_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n284_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G120gat), .B(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT5), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n297_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT13), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT75), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(KEYINPUT75), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n307_), .B2(new_n305_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT76), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G29gat), .B(G36gat), .Z(new_n315_));
  XOR2_X1   g114(.A(G43gat), .B(G50gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT15), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n244_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n317_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n244_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G232gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT34), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT35), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(KEYINPUT35), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT77), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n327_), .B2(KEYINPUT79), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G190gat), .B(G218gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G134gat), .B(G162gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(KEYINPUT36), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(new_n331_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n335_), .B(KEYINPUT36), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT37), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT37), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G15gat), .B(G22gat), .ZN(new_n349_));
  INV_X1    g148(.A(G1gat), .ZN(new_n350_));
  INV_X1    g149(.A(G8gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT14), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G1gat), .B(G8gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G231gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT80), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(new_n267_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n267_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G127gat), .B(G155gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT16), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G183gat), .B(G211gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT17), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n357_), .A2(new_n262_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n364_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n262_), .B2(new_n357_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n348_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n314_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n318_), .A2(new_n355_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n322_), .A2(new_n355_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G229gat), .A2(G233gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n322_), .B(new_n355_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G113gat), .B(G141gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(G169gat), .B(G197gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n383_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT25), .B(G183gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT26), .B(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT83), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT23), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G183gat), .A3(G190gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OR3_X1    g205(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n400_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n399_), .A2(KEYINPUT83), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(KEYINPUT84), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n411_), .B(new_n413_), .C1(KEYINPUT84), .C2(new_n404_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G169gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418_));
  INV_X1    g217(.A(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n410_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(G15gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT30), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n421_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n429_));
  OR3_X1    g228(.A1(new_n423_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n423_), .B2(new_n429_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT85), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G113gat), .B(G120gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT86), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n435_), .A2(KEYINPUT86), .A3(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT31), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n433_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n433_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G22gat), .B(G50gat), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT1), .Z(new_n452_));
  NOR2_X1   g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT88), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n454_), .A2(new_n451_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n456_), .B(KEYINPUT3), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n458_), .B(KEYINPUT2), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(KEYINPUT89), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT89), .B1(new_n461_), .B2(new_n462_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(KEYINPUT89), .A3(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT90), .B1(new_n472_), .B2(new_n460_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n459_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT28), .B1(new_n474_), .B2(KEYINPUT29), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n476_));
  INV_X1    g275(.A(new_n459_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n466_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(KEYINPUT90), .A3(new_n460_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n476_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(new_n475_), .B2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n450_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n449_), .A3(new_n484_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n474_), .A2(KEYINPUT29), .ZN(new_n492_));
  XOR2_X1   g291(.A(G197gat), .B(G204gat), .Z(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT21), .ZN(new_n494_));
  XOR2_X1   g293(.A(G211gat), .B(G218gat), .Z(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n497_));
  INV_X1    g296(.A(G204gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(G197gat), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT21), .B(new_n499_), .C1(new_n493_), .C2(new_n497_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n493_), .A2(KEYINPUT21), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n496_), .A2(new_n500_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n491_), .B1(new_n492_), .B2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n491_), .B(new_n503_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G228gat), .ZN(new_n507_));
  INV_X1    g306(.A(G233gat), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n504_), .A2(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n503_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT92), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n507_), .A2(new_n508_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n505_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n509_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n512_), .A2(new_n513_), .A3(new_n505_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n513_), .B1(new_n512_), .B2(new_n505_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n509_), .A2(KEYINPUT95), .A3(new_n510_), .A4(new_n514_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n490_), .A2(new_n517_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n515_), .A3(KEYINPUT94), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n487_), .A2(new_n489_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n509_), .A2(new_n526_), .A3(new_n510_), .A4(new_n514_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G29gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G85gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT0), .B(G57gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n474_), .A2(new_n536_), .A3(new_n443_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n438_), .A2(new_n440_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n459_), .C1(new_n467_), .C2(new_n473_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n443_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(KEYINPUT4), .C1(new_n544_), .C2(new_n480_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n535_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n545_), .A2(new_n535_), .A3(new_n539_), .A4(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n474_), .A2(new_n443_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n543_), .A3(new_n538_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n534_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n545_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT99), .B1(new_n552_), .B2(new_n540_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n553_), .A2(new_n533_), .A3(new_n549_), .A4(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G226gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT19), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT96), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n502_), .B(new_n417_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n411_), .B(new_n407_), .C1(KEYINPUT84), .C2(new_n404_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n399_), .A2(KEYINPUT98), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n406_), .A2(new_n413_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n416_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n503_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n561_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT97), .B1(new_n560_), .B2(KEYINPUT20), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n559_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n502_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n558_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n563_), .A2(new_n565_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n502_), .B(new_n568_), .C1(new_n577_), .C2(new_n562_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(KEYINPUT20), .A3(new_n576_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G8gat), .B(G36gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT18), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G64gat), .B(G92gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT27), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n560_), .A2(KEYINPUT20), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n559_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n570_), .A4(new_n561_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n578_), .A2(KEYINPUT20), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n558_), .B1(new_n596_), .B2(new_n574_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n584_), .B(KEYINPUT101), .Z(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT27), .B(new_n587_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n529_), .A2(new_n556_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n554_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n545_), .A2(new_n538_), .A3(new_n537_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n548_), .A2(new_n543_), .A3(new_n539_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n534_), .A3(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n586_), .A2(new_n609_), .A3(new_n587_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n547_), .A2(new_n549_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n611_), .A2(KEYINPUT33), .A3(new_n533_), .A4(new_n553_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n606_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n584_), .A2(KEYINPUT32), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT100), .B1(new_n598_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n617_), .B(new_n614_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n618_));
  OAI22_X1  g417(.A1(new_n616_), .A2(new_n618_), .B1(new_n580_), .B2(new_n615_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n554_), .B2(new_n551_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n528_), .B(new_n523_), .C1(new_n613_), .C2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n448_), .B1(new_n604_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n448_), .ZN(new_n623_));
  NOR4_X1   g422(.A1(new_n529_), .A2(new_n555_), .A3(new_n623_), .A4(new_n602_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT102), .B(new_n390_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n624_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(new_n389_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n373_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n350_), .A3(new_n555_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n339_), .A2(KEYINPUT103), .A3(new_n342_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT103), .B1(new_n339_), .B2(new_n342_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n627_), .A2(new_n636_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n389_), .B(new_n371_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n555_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G1gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n629_), .A2(new_n351_), .A3(new_n602_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n637_), .A2(new_n602_), .A3(new_n638_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n648_), .A3(G8gat), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n643_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n643_), .B(KEYINPUT40), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  NAND3_X1  g455(.A1(new_n637_), .A2(new_n448_), .A3(new_n638_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G15gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n629_), .A2(new_n425_), .A3(new_n448_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n629_), .A2(new_n664_), .A3(new_n529_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n637_), .A2(new_n529_), .A3(new_n638_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G22gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1327gat));
  NAND3_X1  g471(.A1(new_n312_), .A2(new_n636_), .A3(new_n371_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n628_), .B2(new_n625_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n556_), .A2(G29gat), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT109), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678_));
  INV_X1    g477(.A(new_n371_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n309_), .A2(new_n389_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n348_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT43), .B1(new_n681_), .B2(new_n682_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n680_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n678_), .B1(new_n689_), .B2(new_n555_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n687_), .A2(new_n678_), .A3(new_n555_), .A4(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n677_), .B1(new_n690_), .B2(new_n692_), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n602_), .A3(new_n688_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n603_), .A2(G36gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n674_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(KEYINPUT46), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n687_), .A2(new_n448_), .A3(new_n688_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G43gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n674_), .A2(new_n419_), .A3(new_n448_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(KEYINPUT47), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  INV_X1    g510(.A(new_n529_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(G50gat), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n674_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n687_), .A2(new_n529_), .A3(new_n688_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G50gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT110), .ZN(G1331gat));
  NOR3_X1   g516(.A1(new_n314_), .A2(new_n390_), .A3(new_n371_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n637_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n556_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n627_), .A2(new_n390_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n312_), .A2(new_n371_), .A3(new_n348_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n253_), .A3(new_n555_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n720_), .A2(new_n725_), .ZN(G1332gat));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n251_), .A3(new_n602_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  INV_X1    g527(.A(new_n719_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n602_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(G64gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT48), .B(new_n251_), .C1(new_n729_), .C2(new_n602_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1333gat));
  OR3_X1    g532(.A1(new_n723_), .A2(G71gat), .A3(new_n623_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n729_), .A2(new_n448_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  NAND3_X1  g538(.A1(new_n724_), .A2(new_n249_), .A3(new_n529_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n729_), .A2(new_n529_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n249_), .C1(new_n729_), .C2(new_n529_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  NOR3_X1   g544(.A1(new_n314_), .A2(new_n679_), .A3(new_n635_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n721_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n555_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n683_), .A2(new_n684_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n390_), .A2(new_n679_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n312_), .A2(KEYINPUT112), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT112), .B1(new_n312_), .B2(new_n755_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n751_), .A2(new_n753_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n555_), .A2(G85gat), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT113), .Z(new_n761_));
  AOI21_X1  g560(.A(new_n749_), .B1(new_n759_), .B2(new_n761_), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n748_), .A2(new_n210_), .A3(new_n602_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n759_), .A2(new_n602_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n210_), .ZN(G1337gat));
  OR2_X1    g564(.A1(new_n623_), .A2(new_n214_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n747_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n751_), .A2(new_n753_), .A3(new_n448_), .A4(new_n758_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G99gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n769_), .B(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n748_), .A2(new_n221_), .A3(new_n529_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n758_), .B(new_n529_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n773_), .B(new_n780_), .C1(new_n777_), .C2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NOR2_X1   g581(.A1(new_n529_), .A2(new_n602_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n623_), .A2(new_n556_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT119), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n374_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n378_), .A2(new_n376_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n386_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n386_), .B2(new_n381_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT117), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n295_), .A2(new_n296_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n302_), .B1(new_n793_), .B2(new_n283_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n284_), .B(new_n301_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT118), .B(new_n792_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n283_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n269_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n244_), .B2(new_n267_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n244_), .A2(new_n275_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n277_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n244_), .A2(KEYINPUT73), .A3(new_n275_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n273_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n283_), .A2(new_n802_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n270_), .B(new_n271_), .C1(new_n276_), .C2(new_n282_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n292_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n803_), .A2(new_n810_), .A3(new_n811_), .A4(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n301_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n301_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT116), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n301_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT116), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n389_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n817_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n635_), .B(new_n787_), .C1(new_n800_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n296_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT72), .B1(new_n291_), .B2(new_n292_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n283_), .B(new_n302_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n827_), .A2(new_n792_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n827_), .B2(new_n792_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n829_), .A2(new_n830_), .B1(new_n816_), .B2(new_n815_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT58), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n833_), .ZN(new_n835_));
  OAI221_X1 g634(.A(new_n835_), .B1(new_n815_), .B2(new_n816_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n348_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n798_), .B(new_n799_), .C1(new_n817_), .C2(new_n822_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n787_), .B1(new_n839_), .B2(new_n635_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n371_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n372_), .A2(new_n842_), .A3(new_n389_), .A4(new_n312_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n347_), .A2(new_n389_), .A3(new_n679_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n309_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n785_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n390_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n846_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n785_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n854_));
  AND4_X1   g653(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .A4(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n851_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(KEYINPUT122), .A3(new_n852_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n847_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(KEYINPUT123), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n390_), .A2(G113gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n848_), .B1(new_n862_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n312_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n847_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n314_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n847_), .B2(new_n679_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n679_), .A2(G127gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n862_), .B2(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n847_), .B2(new_n636_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n348_), .A2(G134gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n862_), .B2(new_n874_), .ZN(G1343gat));
  AOI21_X1  g674(.A(new_n448_), .B1(new_n841_), .B2(new_n846_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n712_), .A2(new_n556_), .A3(new_n602_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n390_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n313_), .A3(new_n311_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n679_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n878_), .A2(new_n886_), .A3(new_n636_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n878_), .A2(new_n348_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n529_), .A2(new_n603_), .A3(new_n623_), .A4(new_n555_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n850_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n389_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT22), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n396_), .B1(new_n893_), .B2(new_n890_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1348gat));
  INV_X1    g697(.A(new_n892_), .ZN(new_n899_));
  AOI21_X1  g698(.A(G176gat), .B1(new_n899_), .B2(new_n309_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n892_), .A2(new_n397_), .A3(new_n314_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n902_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n900_), .B1(new_n903_), .B2(new_n904_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n892_), .A2(new_n371_), .ZN(new_n906_));
  MUX2_X1   g705(.A(G183gat), .B(new_n391_), .S(new_n906_), .Z(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n892_), .B2(new_n347_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n636_), .A2(new_n392_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT125), .Z(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n892_), .B2(new_n910_), .ZN(G1351gat));
  NOR3_X1   g710(.A1(new_n712_), .A2(new_n555_), .A3(new_n603_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n876_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n389_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n314_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n498_), .ZN(G1353gat));
  NOR3_X1   g716(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n918_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n371_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT126), .Z(new_n923_));
  NAND3_X1  g722(.A1(new_n876_), .A2(new_n912_), .A3(new_n923_), .ZN(new_n924_));
  MUX2_X1   g723(.A(new_n918_), .B(new_n921_), .S(new_n924_), .Z(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n913_), .B2(new_n347_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n635_), .A2(G218gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n913_), .B2(new_n927_), .ZN(G1355gat));
endmodule


