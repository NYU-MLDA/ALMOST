//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n970_, new_n972_, new_n973_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1020_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1028_, new_n1029_, new_n1030_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT93), .ZN(new_n203_));
  XOR2_X1   g002(.A(G211gat), .B(G218gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(KEYINPUT91), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT21), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT21), .B2(new_n206_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(KEYINPUT87), .ZN(new_n214_));
  NOR3_X1   g013(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT2), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n218_), .C1(KEYINPUT3), .C2(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(KEYINPUT1), .B2(new_n220_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n213_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n217_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n211_), .B1(new_n231_), .B2(KEYINPUT29), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G228gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT90), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n203_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n208_), .B1(new_n207_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(KEYINPUT21), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n229_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n234_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT93), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(KEYINPUT92), .A3(new_n234_), .A4(new_n240_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n235_), .A2(new_n245_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n250_), .A2(KEYINPUT94), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n235_), .A2(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n249_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT28), .B1(new_n231_), .B2(KEYINPUT29), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n241_), .A2(new_n258_), .A3(new_n242_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G22gat), .B(G50gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n253_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT94), .B1(new_n250_), .B2(new_n252_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n254_), .A2(new_n255_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n251_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n256_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT89), .B1(new_n262_), .B2(new_n263_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n263_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n261_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n266_), .A2(new_n267_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT85), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282_));
  XOR2_X1   g081(.A(G113gat), .B(G120gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT84), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n282_), .A2(new_n283_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n281_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n231_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n284_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n224_), .A2(new_n230_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT96), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT96), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n241_), .A2(new_n297_), .A3(new_n293_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n291_), .A2(new_n295_), .A3(new_n296_), .A4(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G29gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G85gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT0), .B(G57gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n281_), .A2(new_n286_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n292_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n288_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT4), .B1(new_n306_), .B2(new_n231_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n291_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n296_), .B(KEYINPUT97), .Z(new_n310_));
  OAI211_X1 g109(.A(new_n299_), .B(new_n303_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  OR3_X1    g117(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n319_), .A2(KEYINPUT24), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G190gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT95), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT24), .B1(new_n319_), .B2(new_n320_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT23), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n322_), .A2(new_n328_), .A3(KEYINPUT95), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n342_));
  OAI21_X1  g141(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n343_));
  OR3_X1    g142(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n318_), .B1(new_n346_), .B2(new_n240_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n327_), .A2(KEYINPUT81), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(new_n326_), .A3(G190gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n323_), .A2(new_n348_), .A3(new_n325_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n322_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(KEYINPUT83), .A3(new_n322_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n337_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n211_), .A2(new_n345_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n317_), .B1(new_n347_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n240_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n211_), .B1(new_n356_), .B2(new_n345_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n363_), .A3(new_n317_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n360_), .A2(new_n362_), .A3(new_n316_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n358_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n308_), .A2(KEYINPUT4), .ZN(new_n373_));
  INV_X1    g172(.A(new_n307_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n373_), .A2(new_n374_), .B1(G225gat), .B2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n303_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n369_), .B(new_n372_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n313_), .A2(new_n314_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n359_), .A2(new_n364_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n347_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n357_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n316_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n317_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n381_), .B1(new_n386_), .B2(new_n380_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n299_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n376_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n311_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n276_), .B1(new_n379_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT98), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n369_), .A2(KEYINPUT27), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n370_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT99), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(KEYINPUT99), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n369_), .A2(new_n372_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(KEYINPUT27), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n389_), .A2(new_n311_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n268_), .A2(new_n402_), .A3(new_n251_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n267_), .A2(new_n403_), .A3(new_n264_), .A4(new_n256_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n256_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n250_), .A2(new_n252_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n275_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n276_), .B(new_n410_), .C1(new_n379_), .C2(new_n390_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n392_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G43gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT30), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(G15gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n415_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n356_), .A2(new_n345_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT86), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n306_), .B(KEYINPUT31), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n424_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n412_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n397_), .A2(new_n399_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n401_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n404_), .A2(new_n407_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G113gat), .B(G141gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G169gat), .B(G197gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  INV_X1    g240(.A(G36gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G29gat), .ZN(new_n443_));
  INV_X1    g242(.A(G29gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G36gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G43gat), .B(G50gat), .Z(new_n450_));
  NOR3_X1   g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G43gat), .B(G50gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n444_), .A2(G36gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n442_), .A2(G29gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT71), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n455_), .B2(new_n447_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n441_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n450_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n447_), .A3(new_n452_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT15), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT14), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT75), .B(G8gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(G1gat), .ZN(new_n464_));
  INV_X1    g263(.A(G22gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n417_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G15gat), .A2(G22gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT76), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(G1gat), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT14), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n468_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G8gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  AOI221_X4 g278(.A(KEYINPUT76), .B1(new_n466_), .B2(new_n467_), .C1(new_n473_), .C2(KEYINPUT14), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n475_), .B1(new_n474_), .B2(new_n468_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n461_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n470_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n477_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n451_), .A2(new_n456_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT79), .B1(new_n458_), .B2(new_n459_), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n484_), .A2(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n483_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n486_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT79), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n482_), .A2(new_n492_), .A3(new_n478_), .A4(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n440_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n494_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n490_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n482_), .A2(new_n478_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n493_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n483_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n503_), .A3(new_n439_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT80), .Z(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT6), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526_));
  INV_X1    g325(.A(G99gat), .ZN(new_n527_));
  INV_X1    g326(.A(G106gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n530_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n533_), .A2(new_n534_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(KEYINPUT67), .A3(new_n530_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n519_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n532_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n451_), .A2(new_n456_), .ZN(new_n540_));
  OR2_X1    g339(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n528_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT64), .B(G92gat), .ZN(new_n544_));
  INV_X1    g343(.A(G85gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT9), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n543_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n512_), .A2(new_n514_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n525_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT65), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n516_), .A2(new_n517_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n553_), .A2(KEYINPUT9), .B1(new_n522_), .B2(new_n524_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT64), .B(G92gat), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n546_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT65), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .A4(new_n543_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n539_), .A2(new_n540_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n509_), .A2(new_n510_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n539_), .A2(new_n559_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n511_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT73), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n566_), .B(KEYINPUT72), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n565_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n539_), .A2(new_n559_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n461_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n511_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n561_), .A4(new_n560_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n564_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n564_), .A2(new_n582_), .A3(KEYINPUT74), .A4(new_n578_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n576_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(KEYINPUT36), .A3(new_n574_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n577_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n564_), .B2(new_n582_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n530_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n534_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n525_), .A3(new_n536_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n519_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n603_), .A2(KEYINPUT8), .B1(new_n531_), .B2(new_n520_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n552_), .A2(new_n558_), .ZN(new_n605_));
  INV_X1    g404(.A(G71gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G78gat), .ZN(new_n607_));
  INV_X1    g406(.A(G78gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G71gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G57gat), .B(G64gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(KEYINPUT11), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT68), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n611_), .B2(KEYINPUT11), .ZN(new_n614_));
  INV_X1    g413(.A(G64gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G57gat), .ZN(new_n616_));
  INV_X1    g415(.A(G57gat), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G64gat), .ZN(new_n618_));
  AND4_X1   g417(.A1(new_n613_), .A2(new_n616_), .A3(new_n618_), .A4(KEYINPUT11), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n612_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n618_), .A3(KEYINPUT11), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT68), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n618_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT11), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n616_), .A2(new_n618_), .A3(new_n613_), .A4(KEYINPUT11), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n622_), .A2(new_n625_), .A3(new_n610_), .A4(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n620_), .A2(new_n627_), .A3(KEYINPUT69), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT69), .B1(new_n620_), .B2(new_n627_), .ZN(new_n629_));
  OAI22_X1  g428(.A1(new_n604_), .A2(new_n605_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n603_), .A2(KEYINPUT8), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n635_), .A2(new_n532_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n628_), .A2(new_n629_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n620_), .A2(new_n627_), .A3(KEYINPUT12), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n539_), .B2(new_n559_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n638_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n620_), .A2(new_n627_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT69), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n620_), .A2(new_n627_), .A3(KEYINPUT69), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n579_), .A2(new_n647_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n559_), .A2(new_n539_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n634_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT5), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n652_), .B(new_n653_), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n642_), .A2(new_n650_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n642_), .B2(new_n650_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n597_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n642_), .A2(new_n650_), .A3(new_n655_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT13), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT70), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(G127gat), .B(G155gat), .Z(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G183gat), .B(G211gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT17), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT78), .ZN(new_n672_));
  INV_X1    g471(.A(new_n500_), .ZN(new_n673_));
  AND2_X1   g472(.A1(G231gat), .A2(G233gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n674_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n647_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n637_), .B1(new_n679_), .B2(new_n675_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n643_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n679_), .B2(new_n675_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(new_n677_), .A3(new_n643_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(KEYINPUT17), .A4(new_n669_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n591_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT37), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n595_), .A2(new_n664_), .A3(new_n687_), .A4(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n436_), .A2(new_n506_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G1gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n401_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n202_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT102), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n434_), .B1(new_n412_), .B2(new_n428_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n506_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n690_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(KEYINPUT38), .A3(new_n693_), .A4(new_n401_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n664_), .A2(new_n505_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n686_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n401_), .B(new_n381_), .C1(new_n386_), .C2(new_n380_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n311_), .A2(new_n312_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n311_), .A2(new_n312_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n375_), .A2(new_n377_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n398_), .A4(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n433_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n710_), .A2(new_n410_), .B1(new_n400_), .B2(new_n408_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n427_), .B1(new_n711_), .B2(new_n392_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n593_), .B(new_n704_), .C1(new_n712_), .C2(new_n434_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G1gat), .B1(new_n713_), .B2(new_n431_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n696_), .A2(new_n702_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n696_), .A2(new_n702_), .A3(KEYINPUT103), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1324gat));
  OR3_X1    g520(.A1(new_n692_), .A2(new_n400_), .A3(new_n463_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT39), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n697_), .A2(new_n688_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n724_), .A2(KEYINPUT104), .A3(new_n430_), .A4(new_n704_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(G8gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n713_), .B2(new_n400_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n723_), .A2(new_n728_), .A3(new_n725_), .A4(G8gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n722_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT40), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT40), .B(new_n722_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1325gat));
  OAI21_X1  g534(.A(G15gat), .B1(new_n713_), .B2(new_n428_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT41), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n699_), .A2(new_n417_), .A3(new_n427_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1326gat));
  OAI21_X1  g538(.A(G22gat), .B1(new_n713_), .B2(new_n276_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT42), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n699_), .A2(new_n465_), .A3(new_n433_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1327gat));
  NOR2_X1   g542(.A1(new_n697_), .A2(new_n698_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n664_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n686_), .A2(new_n688_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G29gat), .B1(new_n749_), .B2(new_n401_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT37), .B1(new_n587_), .B2(new_n592_), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n594_), .B(new_n591_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n697_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n755_));
  INV_X1    g554(.A(new_n753_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n755_), .B(new_n756_), .C1(new_n712_), .C2(new_n434_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n703_), .A2(new_n687_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT44), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n761_));
  INV_X1    g560(.A(new_n759_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n761_), .B(new_n762_), .C1(new_n754_), .C2(new_n757_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n431_), .A2(new_n444_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n750_), .B1(new_n764_), .B2(new_n765_), .ZN(G1328gat));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n442_), .B1(new_n764_), .B2(new_n430_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n400_), .A2(G36gat), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n748_), .A2(KEYINPUT45), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT45), .B1(new_n748_), .B2(new_n770_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n768_), .B2(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n760_), .A2(new_n763_), .A3(new_n400_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT46), .B(new_n773_), .C1(new_n776_), .C2(new_n442_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1329gat));
  INV_X1    g577(.A(G43gat), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n428_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n764_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n748_), .B2(new_n428_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT47), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1330gat));
  NAND2_X1  g586(.A1(new_n764_), .A2(new_n433_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G50gat), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n276_), .A2(G50gat), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT105), .Z(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n748_), .B2(new_n791_), .ZN(G1331gat));
  NOR2_X1   g591(.A1(new_n697_), .A2(new_n505_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n751_), .A2(new_n752_), .A3(new_n686_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n745_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n796_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n617_), .A3(new_n401_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n506_), .A2(new_n664_), .A3(new_n686_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n436_), .A2(new_n593_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G57gat), .B1(new_n802_), .B2(new_n431_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(G1332gat));
  NAND4_X1  g603(.A1(new_n797_), .A2(new_n798_), .A3(new_n615_), .A4(new_n430_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G64gat), .B1(new_n802_), .B2(new_n400_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT48), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n806_), .A2(KEYINPUT48), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT107), .B(new_n805_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1333gat));
  NAND3_X1  g613(.A1(new_n799_), .A2(new_n606_), .A3(new_n427_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G71gat), .B1(new_n802_), .B2(new_n428_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT49), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1334gat));
  NAND3_X1  g617(.A1(new_n799_), .A2(new_n608_), .A3(new_n433_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G78gat), .B1(new_n802_), .B2(new_n276_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT50), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n746_), .A2(new_n664_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n793_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n545_), .A3(new_n401_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n664_), .A2(new_n687_), .A3(new_n505_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT109), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n758_), .A2(KEYINPUT108), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n754_), .A2(new_n831_), .A3(new_n757_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n401_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n826_), .B1(new_n834_), .B2(new_n545_), .ZN(G1336gat));
  AOI21_X1  g634(.A(G92gat), .B1(new_n825_), .B2(new_n430_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n400_), .A2(new_n544_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n833_), .B2(new_n837_), .ZN(G1337gat));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n427_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n428_), .B(new_n829_), .C1(new_n830_), .C2(new_n832_), .ZN(new_n841_));
  OAI221_X1 g640(.A(new_n839_), .B1(new_n824_), .B2(new_n840_), .C1(new_n841_), .C2(new_n527_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n527_), .B1(new_n833_), .B2(new_n427_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n824_), .A2(new_n840_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(G1338gat));
  NAND3_X1  g645(.A1(new_n825_), .A2(new_n528_), .A3(new_n433_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n829_), .A2(new_n276_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n528_), .B1(new_n758_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT53), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n847_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1339gat));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n690_), .B2(new_n506_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n794_), .A2(new_n859_), .A3(new_n664_), .A4(new_n698_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n640_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n648_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n633_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n642_), .A2(KEYINPUT55), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n867_), .A3(new_n638_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n865_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n869_), .B2(new_n655_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT111), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n655_), .A2(new_n862_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n869_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n863_), .A2(new_n864_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n634_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n868_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n867_), .B1(new_n863_), .B2(new_n638_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT111), .A3(new_n872_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n870_), .A2(new_n874_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n505_), .A2(new_n660_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT110), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n884_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n497_), .A2(new_n498_), .B1(new_n502_), .B2(new_n483_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n439_), .B1(new_n497_), .B2(new_n490_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n483_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n886_), .A2(new_n439_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT112), .B(new_n889_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(KEYINPUT57), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n593_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n894_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(new_n688_), .ZN(new_n902_));
  AND4_X1   g701(.A1(new_n478_), .A2(new_n482_), .A3(new_n493_), .A4(new_n492_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n482_), .A2(new_n478_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n490_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n440_), .A3(new_n888_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n504_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT114), .B1(new_n656_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n889_), .A2(new_n909_), .A3(new_n660_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n879_), .A2(new_n872_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n870_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n914_), .A3(KEYINPUT58), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n917_), .A2(new_n756_), .A3(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n900_), .A2(new_n902_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n861_), .B1(new_n920_), .B2(new_n686_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR4_X1   g721(.A1(new_n430_), .A2(new_n433_), .A3(new_n431_), .A4(new_n428_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT115), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n922_), .A2(new_n926_), .A3(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(G113gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n505_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n924_), .B1(KEYINPUT116), .B2(KEYINPUT59), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(KEYINPUT116), .B2(KEYINPUT59), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n924_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n698_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n931_), .B1(new_n937_), .B2(new_n930_), .ZN(G1340gat));
  INV_X1    g737(.A(G120gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n929_), .B(new_n940_), .C1(KEYINPUT60), .C2(new_n939_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n664_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n939_), .ZN(G1341gat));
  INV_X1    g742(.A(G127gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n928_), .B2(new_n686_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT117), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  OAI211_X1 g746(.A(KEYINPUT117), .B(new_n944_), .C1(new_n928_), .C2(new_n686_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n933_), .A2(new_n936_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT118), .B(G127gat), .Z(new_n950_));
  AND2_X1   g749(.A1(new_n687_), .A2(new_n950_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n947_), .A2(new_n948_), .B1(new_n949_), .B2(new_n951_), .ZN(G1342gat));
  AOI21_X1  g751(.A(G134gat), .B1(new_n929_), .B2(new_n688_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n756_), .A2(G134gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT119), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n949_), .B2(new_n955_), .ZN(G1343gat));
  NAND4_X1  g755(.A1(new_n400_), .A2(new_n401_), .A3(new_n433_), .A4(new_n428_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT120), .B1(new_n921_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n959_));
  INV_X1    g758(.A(new_n957_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n688_), .B1(new_n885_), .B2(new_n895_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n911_), .B1(new_n913_), .B2(new_n870_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n753_), .B1(new_n962_), .B2(KEYINPUT58), .ZN(new_n963_));
  AOI22_X1  g762(.A1(new_n961_), .A2(new_n899_), .B1(new_n963_), .B2(new_n917_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n687_), .B1(new_n964_), .B2(new_n902_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n959_), .B(new_n960_), .C1(new_n965_), .C2(new_n861_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n958_), .A2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(new_n505_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n745_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g770(.A1(new_n967_), .A2(new_n687_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(KEYINPUT61), .B(G155gat), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n972_), .B(new_n973_), .ZN(G1346gat));
  NAND3_X1  g773(.A1(new_n967_), .A2(G162gat), .A3(new_n756_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n967_), .A2(new_n688_), .ZN(new_n977_));
  INV_X1    g776(.A(G162gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n976_), .B1(new_n977_), .B2(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n593_), .B1(new_n958_), .B2(new_n966_), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n980_), .A2(KEYINPUT121), .A3(G162gat), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n975_), .B1(new_n979_), .B2(new_n981_), .ZN(new_n982_));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  OAI211_X1 g783(.A(KEYINPUT122), .B(new_n975_), .C1(new_n979_), .C2(new_n981_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(G1347gat));
  NOR4_X1   g785(.A1(new_n921_), .A2(new_n433_), .A3(new_n400_), .A4(new_n432_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n987_), .A2(new_n505_), .ZN(new_n988_));
  XOR2_X1   g787(.A(KEYINPUT22), .B(G169gat), .Z(new_n989_));
  NOR2_X1   g788(.A1(new_n988_), .A2(new_n989_), .ZN(new_n990_));
  AOI21_X1  g789(.A(KEYINPUT123), .B1(new_n988_), .B2(G169gat), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n990_), .B1(new_n991_), .B2(new_n992_), .ZN(new_n993_));
  OR2_X1    g792(.A1(new_n991_), .A2(new_n992_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n988_), .A2(G169gat), .ZN(new_n995_));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n996_));
  NOR2_X1   g795(.A1(new_n995_), .A2(new_n996_), .ZN(new_n997_));
  OAI21_X1  g796(.A(new_n993_), .B1(new_n994_), .B2(new_n997_), .ZN(G1348gat));
  XNOR2_X1  g797(.A(KEYINPUT124), .B(G176gat), .ZN(new_n999_));
  INV_X1    g798(.A(G176gat), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(new_n1000_), .A2(KEYINPUT124), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n987_), .A2(new_n745_), .ZN(new_n1002_));
  MUX2_X1   g801(.A(new_n999_), .B(new_n1001_), .S(new_n1002_), .Z(G1349gat));
  NAND2_X1  g802(.A1(new_n987_), .A2(new_n687_), .ZN(new_n1004_));
  INV_X1    g803(.A(G183gat), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1004_), .A2(new_n1005_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1006_), .B1(new_n323_), .B2(new_n1004_), .ZN(new_n1007_));
  XNOR2_X1  g806(.A(new_n1007_), .B(KEYINPUT125), .ZN(G1350gat));
  NAND4_X1  g807(.A1(new_n987_), .A2(new_n325_), .A3(new_n327_), .A4(new_n688_), .ZN(new_n1009_));
  AND2_X1   g808(.A1(new_n987_), .A2(new_n756_), .ZN(new_n1010_));
  OAI21_X1  g809(.A(new_n1009_), .B1(new_n1010_), .B2(new_n324_), .ZN(G1351gat));
  AND3_X1   g810(.A1(new_n430_), .A2(new_n408_), .A3(new_n428_), .ZN(new_n1012_));
  AND2_X1   g811(.A1(new_n922_), .A2(new_n1012_), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(new_n1013_), .A2(new_n505_), .ZN(new_n1014_));
  INV_X1    g813(.A(G197gat), .ZN(new_n1015_));
  NOR3_X1   g814(.A1(new_n1014_), .A2(KEYINPUT126), .A3(new_n1015_), .ZN(new_n1016_));
  NAND3_X1  g815(.A1(new_n1013_), .A2(G197gat), .A3(new_n505_), .ZN(new_n1017_));
  AND2_X1   g816(.A1(new_n1017_), .A2(KEYINPUT126), .ZN(new_n1018_));
  AOI211_X1 g817(.A(new_n1016_), .B(new_n1018_), .C1(new_n1015_), .C2(new_n1014_), .ZN(G1352gat));
  NAND2_X1  g818(.A1(new_n1013_), .A2(new_n745_), .ZN(new_n1020_));
  XNOR2_X1  g819(.A(new_n1020_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g820(.A1(new_n922_), .A2(new_n687_), .A3(new_n1012_), .ZN(new_n1022_));
  NOR3_X1   g821(.A1(new_n1022_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023_));
  OR2_X1    g822(.A1(new_n1023_), .A2(KEYINPUT127), .ZN(new_n1024_));
  NAND2_X1  g823(.A1(new_n1023_), .A2(KEYINPUT127), .ZN(new_n1025_));
  XOR2_X1   g824(.A(KEYINPUT63), .B(G211gat), .Z(new_n1026_));
  AOI22_X1  g825(.A1(new_n1024_), .A2(new_n1025_), .B1(new_n1022_), .B2(new_n1026_), .ZN(G1354gat));
  INV_X1    g826(.A(G218gat), .ZN(new_n1028_));
  NAND3_X1  g827(.A1(new_n1013_), .A2(new_n1028_), .A3(new_n688_), .ZN(new_n1029_));
  AND2_X1   g828(.A1(new_n1013_), .A2(new_n756_), .ZN(new_n1030_));
  OAI21_X1  g829(.A(new_n1029_), .B1(new_n1030_), .B2(new_n1028_), .ZN(G1355gat));
endmodule


