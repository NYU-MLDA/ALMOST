//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G85gat), .B(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT67), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(KEYINPUT67), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  MUX2_X1   g019(.A(KEYINPUT9), .B(new_n220_), .S(new_n208_), .Z(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n204_), .A3(new_n224_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT71), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(KEYINPUT15), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT34), .Z(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G190gat), .B(G218gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT73), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G134gat), .B(G162gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT36), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT74), .Z(new_n250_));
  NOR2_X1   g049(.A1(new_n239_), .A2(new_n240_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n237_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT72), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(KEYINPUT72), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n243_), .B(new_n250_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT75), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n202_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n255_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n242_), .B1(new_n259_), .B2(new_n253_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n247_), .B(new_n248_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  OAI221_X1 g062(.A(new_n256_), .B1(new_n257_), .B2(new_n202_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT76), .B(G1gat), .ZN(new_n266_));
  INV_X1    g065(.A(G8gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G15gat), .B(G22gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT77), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G1gat), .B(G8gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n270_), .B(KEYINPUT77), .ZN(new_n275_));
  INV_X1    g074(.A(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n281_));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n278_), .B(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G127gat), .B(G155gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT16), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G183gat), .B(G211gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n288_), .A2(new_n294_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n265_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT78), .Z(new_n300_));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT87), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n303_), .B(new_n304_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  AND2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT1), .ZN(new_n313_));
  INV_X1    g112(.A(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n310_), .B1(new_n313_), .B2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n318_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n324_), .A2(new_n327_), .A3(KEYINPUT88), .A4(new_n317_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n314_), .A2(new_n315_), .A3(KEYINPUT89), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT3), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n318_), .A2(KEYINPUT90), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT2), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n318_), .A2(KEYINPUT90), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(KEYINPUT89), .A3(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n333_), .A3(new_n335_), .A4(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n311_), .A2(new_n312_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n309_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n329_), .A2(new_n340_), .A3(new_n307_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n303_), .A2(new_n304_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n303_), .A2(new_n304_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n308_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n305_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n320_), .A2(new_n328_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n344_), .B(KEYINPUT96), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n309_), .A2(new_n341_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT97), .B1(new_n353_), .B2(KEYINPUT4), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  AOI211_X1 g154(.A(new_n355_), .B(new_n342_), .C1(new_n350_), .C2(new_n352_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n302_), .B(new_n343_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  AOI21_X1  g160(.A(new_n302_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT98), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n357_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n357_), .B2(new_n363_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n236_), .A2(new_n278_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G229gat), .A2(G233gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n278_), .A2(new_n234_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(KEYINPUT79), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n274_), .A2(new_n277_), .A3(new_n233_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT80), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n378_), .A3(new_n375_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n371_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G141gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G169gat), .B(G197gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  AND2_X1   g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n380_), .A2(new_n383_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT81), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT26), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT82), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n393_), .A4(new_n389_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT23), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n408_), .B(new_n412_), .C1(KEYINPUT24), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G183gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n395_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n406_), .A2(new_n419_), .A3(new_n407_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G169gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n408_), .A2(KEYINPUT84), .A3(new_n419_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n403_), .A2(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT30), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT86), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT85), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(new_n309_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n428_), .A2(KEYINPUT86), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT31), .Z(new_n439_));
  OR2_X1    g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n439_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n367_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(G197gat), .A2(G204gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT21), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(KEYINPUT21), .A3(new_n446_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G211gat), .B(G218gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n450_), .A2(new_n451_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n341_), .B2(KEYINPUT29), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G78gat), .B(G106gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n341_), .A2(KEYINPUT29), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT28), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n463_), .B(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n460_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n427_), .B2(new_n455_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n411_), .B(KEYINPUT93), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n413_), .A2(KEYINPUT22), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT22), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G169gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n420_), .B(new_n476_), .C1(new_n483_), .C2(G176gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT26), .B(G190gat), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n485_), .A2(new_n389_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n406_), .A2(new_n407_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n415_), .A2(KEYINPUT24), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n484_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n454_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n473_), .B1(new_n475_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n416_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n426_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n454_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n455_), .B(new_n484_), .C1(new_n488_), .C2(new_n492_), .ZN(new_n499_));
  AND4_X1   g298(.A1(KEYINPUT20), .A2(new_n498_), .A3(new_n499_), .A4(new_n473_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G8gat), .B(G36gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G64gat), .B(G92gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n470_), .B1(new_n501_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT20), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n472_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n475_), .A2(new_n473_), .A3(new_n494_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT101), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(KEYINPUT101), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n495_), .B2(new_n500_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n403_), .A2(new_n417_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n425_), .A2(new_n426_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n455_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n494_), .A2(new_n520_), .A3(KEYINPUT20), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n472_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT20), .A4(new_n473_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n507_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n517_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n470_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n515_), .A2(new_n516_), .A3(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n444_), .A2(new_n469_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n469_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n357_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n301_), .B(new_n343_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n361_), .B1(new_n353_), .B2(new_n302_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n525_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n357_), .A2(new_n363_), .A3(KEYINPUT33), .A4(new_n361_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n510_), .A2(new_n511_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n507_), .A2(KEYINPUT32), .ZN(new_n539_));
  MUX2_X1   g338(.A(new_n538_), .B(new_n501_), .S(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n357_), .A2(new_n363_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n361_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(new_n530_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n544_), .B2(KEYINPUT99), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n539_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n501_), .B2(new_n539_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT99), .B(new_n547_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n529_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n547_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n548_), .A3(new_n537_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(KEYINPUT100), .A3(new_n529_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n527_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n469_), .A3(new_n366_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n528_), .B1(new_n560_), .B2(new_n442_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT13), .ZN(new_n562_));
  XOR2_X1   g361(.A(G120gat), .B(G148gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n285_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n229_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n229_), .A2(new_n568_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n570_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n573_), .A2(KEYINPUT68), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(KEYINPUT68), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n571_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n581_), .B2(new_n569_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n567_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n582_), .A3(new_n567_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n562_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n583_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n388_), .A2(new_n561_), .A3(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n300_), .A2(new_n266_), .A3(new_n367_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n262_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n561_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n586_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n588_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n380_), .B(new_n383_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n595_), .A2(new_n298_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n366_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n592_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n601_), .A3(new_n602_), .ZN(G1324gat));
  OAI21_X1  g402(.A(G8gat), .B1(new_n600_), .B2(new_n558_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n300_), .A2(new_n590_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n527_), .A2(new_n267_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n606_), .A2(KEYINPUT39), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n604_), .A2(new_n605_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n600_), .B2(new_n442_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n607_), .A2(G15gat), .A3(new_n442_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  XOR2_X1   g417(.A(new_n469_), .B(KEYINPUT104), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G22gat), .B1(new_n600_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(G22gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT106), .Z(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(new_n607_), .B2(new_n625_), .ZN(G1327gat));
  INV_X1    g425(.A(new_n528_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n556_), .A2(KEYINPUT100), .A3(new_n529_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT100), .B1(new_n556_), .B2(new_n529_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n529_), .A2(new_n527_), .A3(new_n367_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n442_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n262_), .A2(new_n298_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(new_n598_), .A3(new_n387_), .A4(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n367_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(new_n298_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n598_), .A2(new_n639_), .A3(new_n599_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT43), .B1(new_n561_), .B2(new_n265_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  INV_X1    g441(.A(new_n265_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n629_), .A2(new_n630_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n632_), .B1(new_n644_), .B2(new_n557_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n642_), .B(new_n643_), .C1(new_n645_), .C2(new_n528_), .ZN(new_n646_));
  AOI211_X1 g445(.A(new_n638_), .B(new_n640_), .C1(new_n641_), .C2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n646_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n640_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n367_), .A2(G29gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n637_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n558_), .A2(G36gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n636_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n635_), .A2(KEYINPUT45), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n642_), .B1(new_n633_), .B2(new_n643_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n561_), .A2(KEYINPUT43), .A3(new_n265_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n649_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n638_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n527_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n660_), .B1(new_n666_), .B2(G36gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n654_), .B1(new_n667_), .B2(KEYINPUT46), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n667_), .B2(KEYINPUT107), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n671_), .B(new_n660_), .C1(new_n666_), .C2(G36gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n651_), .B2(new_n527_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n675_), .B2(new_n660_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n667_), .A2(KEYINPUT107), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n654_), .A4(new_n669_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n673_), .A2(new_n678_), .ZN(G1329gat));
  AOI21_X1  g478(.A(G43gat), .B1(new_n636_), .B2(new_n632_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n632_), .A2(G43gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n651_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(G1330gat));
  AOI21_X1  g483(.A(G50gat), .B1(new_n636_), .B2(new_n619_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n469_), .A2(G50gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n651_), .B2(new_n686_), .ZN(G1331gat));
  NOR3_X1   g486(.A1(new_n561_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n300_), .A2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT110), .Z(new_n690_));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n367_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n595_), .A2(new_n298_), .A3(new_n589_), .A4(new_n388_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n366_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n696_), .A3(new_n527_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G64gat), .B1(new_n693_), .B2(new_n558_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1333gat));
  INV_X1    g500(.A(G71gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n690_), .A2(new_n702_), .A3(new_n632_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G71gat), .B1(new_n693_), .B2(new_n442_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n690_), .A2(new_n708_), .A3(new_n619_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G78gat), .B1(new_n693_), .B2(new_n620_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT50), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n598_), .A2(new_n298_), .A3(new_n599_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n648_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n366_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n688_), .A2(new_n634_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n366_), .A2(G85gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(G1336gat));
  OAI21_X1  g517(.A(new_n219_), .B1(new_n716_), .B2(new_n558_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT113), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n714_), .A2(new_n219_), .A3(new_n558_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1337gat));
  NOR3_X1   g521(.A1(new_n716_), .A2(new_n226_), .A3(new_n442_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT115), .ZN(new_n724_));
  INV_X1    g523(.A(new_n714_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n632_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT114), .B1(new_n726_), .B2(G99gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT116), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n729_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1338gat));
  NOR3_X1   g534(.A1(new_n716_), .A2(G106gat), .A3(new_n529_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT117), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n725_), .A2(new_n469_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G106gat), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g543(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n380_), .A2(new_n383_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n374_), .A2(new_n369_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n369_), .B1(new_n278_), .B2(new_n234_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n383_), .B1(new_n368_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n585_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT120), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n567_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(new_n579_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n576_), .A2(new_n755_), .A3(new_n578_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n745_), .B1(new_n753_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n751_), .B(KEYINPUT120), .ZN(new_n766_));
  INV_X1    g565(.A(new_n745_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n768_), .A3(new_n643_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n386_), .B2(new_n587_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n760_), .B2(KEYINPUT119), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n759_), .A2(new_n774_), .A3(KEYINPUT56), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n599_), .A2(KEYINPUT118), .A3(new_n585_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n771_), .A2(new_n773_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n746_), .B(new_n750_), .C1(new_n587_), .C2(new_n583_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n594_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n769_), .B1(new_n779_), .B2(KEYINPUT57), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(KEYINPUT57), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n639_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n387_), .A2(new_n299_), .A3(new_n589_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT54), .Z(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NOR4_X1   g584(.A1(new_n442_), .A2(new_n527_), .A3(new_n469_), .A4(new_n366_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n599_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(KEYINPUT59), .A3(new_n786_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n388_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(new_n789_), .ZN(G1340gat));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n788_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n796_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n598_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n796_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n788_), .A2(new_n801_), .A3(new_n298_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n639_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1342gat));
  INV_X1    g603(.A(G134gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n788_), .A2(new_n805_), .A3(new_n594_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n265_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n805_), .ZN(G1343gat));
  NOR2_X1   g607(.A1(new_n632_), .A2(new_n529_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n810_), .A2(new_n366_), .A3(new_n527_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n599_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n589_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT123), .B(G148gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NAND3_X1  g617(.A1(new_n785_), .A2(new_n298_), .A3(new_n811_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT124), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n821_), .A3(new_n298_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1346gat));
  INV_X1    g625(.A(new_n813_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n827_), .A2(G162gat), .A3(new_n262_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G162gat), .B1(new_n827_), .B2(new_n265_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1347gat));
  NOR2_X1   g629(.A1(new_n444_), .A2(new_n558_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n599_), .A3(new_n620_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n835_), .A3(G169gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n834_), .A2(new_n483_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n834_), .B2(G169gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1348gat));
  AND2_X1   g638(.A1(new_n833_), .A2(new_n529_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n598_), .A2(new_n414_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n833_), .A2(new_n589_), .A3(new_n620_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n840_), .A2(new_n841_), .B1(new_n842_), .B2(new_n414_), .ZN(G1349gat));
  NAND2_X1  g642(.A1(new_n833_), .A2(new_n620_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(new_n639_), .A3(new_n389_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n833_), .A2(KEYINPUT125), .A3(new_n298_), .A4(new_n529_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(new_n418_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n298_), .A3(new_n529_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n847_), .B2(new_n850_), .ZN(G1350gat));
  OAI21_X1  g650(.A(G190gat), .B1(new_n844_), .B2(new_n265_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n594_), .A2(new_n485_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n844_), .B2(new_n853_), .ZN(G1351gat));
  NOR3_X1   g653(.A1(new_n810_), .A2(new_n367_), .A3(new_n558_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n599_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n589_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n860_), .B(new_n861_), .Z(G1353gat));
  AOI211_X1 g661(.A(KEYINPUT63), .B(G211gat), .C1(new_n857_), .C2(new_n298_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n857_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n639_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT63), .B(G211gat), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n865_), .B2(new_n866_), .ZN(G1354gat));
  INV_X1    g666(.A(KEYINPUT127), .ZN(new_n868_));
  INV_X1    g667(.A(G218gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n857_), .A2(new_n869_), .A3(new_n594_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n857_), .B2(new_n643_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT127), .A3(new_n870_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1355gat));
endmodule


