//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT91), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G197gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT87), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT85), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT21), .B1(new_n209_), .B2(KEYINPUT85), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n205_), .B1(new_n212_), .B2(KEYINPUT21), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT86), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G218gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G211gat), .ZN(new_n225_));
  INV_X1    g024(.A(G211gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G218gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n206_), .B2(new_n214_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT85), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n210_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT21), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n218_), .B1(new_n223_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G183gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT25), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G183gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT26), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n241_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT77), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G169gat), .B2(G176gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT24), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT93), .B1(new_n248_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(new_n250_), .B2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT23), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(G183gat), .A3(G190gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n257_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n238_), .A2(G183gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n236_), .A2(KEYINPUT25), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT92), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n254_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n256_), .A2(new_n262_), .A3(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT78), .B(G176gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT22), .B(G169gat), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n272_), .A2(new_n273_), .B1(G169gat), .B2(G176gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n260_), .B2(new_n258_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n260_), .B2(new_n258_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n235_), .B1(new_n271_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n229_), .A2(new_n233_), .A3(new_n232_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n233_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n217_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n244_), .A2(new_n246_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n254_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n262_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n204_), .B1(new_n279_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT94), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n262_), .A2(new_n284_), .B1(new_n277_), .B2(new_n274_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT95), .B1(new_n235_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n282_), .A2(new_n293_), .A3(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n203_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n271_), .A2(new_n235_), .A3(new_n278_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n295_), .A2(KEYINPUT20), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT94), .B(new_n204_), .C1(new_n279_), .C2(new_n287_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n290_), .A2(new_n304_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT27), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT103), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n279_), .A2(new_n287_), .A3(new_n204_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n313_));
  INV_X1    g112(.A(new_n278_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n270_), .A2(new_n262_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n256_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n316_), .B2(new_n235_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n296_), .B1(new_n317_), .B2(new_n295_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT99), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n312_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT99), .B(new_n296_), .C1(new_n317_), .C2(new_n295_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n310_), .B(new_n305_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n292_), .A2(new_n294_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n297_), .A2(KEYINPUT20), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n203_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n311_), .B1(new_n325_), .B2(KEYINPUT99), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n318_), .A2(new_n319_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n304_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n307_), .A2(new_n310_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n322_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n309_), .B1(new_n330_), .B2(KEYINPUT27), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(new_n342_), .C2(new_n336_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(KEYINPUT83), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n335_), .A2(new_n346_), .A3(new_n336_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n349_));
  NOR4_X1   g148(.A1(new_n349_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT80), .B1(new_n339_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n341_), .A2(KEYINPUT81), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT81), .B1(new_n341_), .B2(new_n353_), .ZN(new_n355_));
  OAI22_X1  g154(.A1(new_n350_), .A2(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT82), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT82), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n348_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n348_), .B(KEYINPUT84), .C1(new_n356_), .C2(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n344_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n282_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n282_), .B2(KEYINPUT88), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  OAI221_X1 g171(.A(new_n282_), .B1(KEYINPUT88), .B2(new_n370_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n334_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n374_), .A2(KEYINPUT89), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n334_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n374_), .B2(KEYINPUT89), .ZN(new_n377_));
  INV_X1    g176(.A(new_n344_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n366_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n380_));
  INV_X1    g179(.A(G141gat), .ZN(new_n381_));
  INV_X1    g180(.A(G148gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n351_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n349_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n339_), .A2(KEYINPUT80), .A3(new_n351_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n341_), .A2(new_n353_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n341_), .A2(KEYINPUT81), .A3(new_n353_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT84), .B1(new_n392_), .B2(new_n348_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n378_), .B1(new_n379_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT28), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n367_), .A2(new_n396_), .A3(new_n368_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n395_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n400_));
  OAI22_X1  g199(.A1(new_n375_), .A2(new_n377_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n374_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n399_), .A2(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n374_), .A2(new_n402_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n376_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n332_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT0), .B(G57gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n378_), .B(new_n418_), .C1(new_n379_), .C2(new_n393_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n418_), .B(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n419_), .B(KEYINPUT4), .C1(new_n367_), .C2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n365_), .A2(new_n366_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n424_), .B2(new_n378_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n418_), .B(KEYINPUT79), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n394_), .A2(new_n423_), .A3(new_n429_), .A4(new_n427_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n415_), .B(new_n422_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n419_), .B(new_n414_), .C1(new_n367_), .C2(new_n421_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n413_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n422_), .A2(new_n415_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n394_), .A2(new_n429_), .A3(new_n427_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT97), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n437_), .B2(new_n430_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n413_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT101), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n422_), .A2(new_n415_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n430_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT101), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n434_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(G15gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT30), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n291_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n429_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  INV_X1    g251(.A(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n446_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n409_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT102), .ZN(new_n460_));
  INV_X1    g259(.A(new_n439_), .ZN(new_n461_));
  OR2_X1    g260(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n432_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n419_), .B(new_n415_), .C1(new_n367_), .C2(new_n421_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n413_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n428_), .A2(new_n431_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n422_), .A2(new_n414_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n443_), .A2(new_n462_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n308_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT100), .B(new_n473_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT100), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n325_), .A2(KEYINPUT99), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n327_), .A3(new_n312_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n473_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n300_), .A2(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n440_), .A2(new_n445_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n433_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n465_), .B1(new_n438_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n481_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n472_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n460_), .B1(new_n486_), .B2(new_n407_), .ZN(new_n487_));
  AOI211_X1 g286(.A(KEYINPUT101), .B(new_n439_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n444_), .B1(new_n432_), .B2(new_n461_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n484_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n478_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT100), .ZN(new_n492_));
  INV_X1    g291(.A(new_n481_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n477_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n470_), .A2(new_n471_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n308_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(KEYINPUT102), .A3(new_n408_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n407_), .A2(new_n446_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT104), .B1(new_n331_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n490_), .B1(new_n401_), .B2(new_n406_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT104), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT27), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n305_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n307_), .A2(new_n310_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n508_), .B2(new_n322_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n503_), .B(new_n504_), .C1(new_n509_), .C2(new_n309_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n487_), .A2(new_n500_), .A3(new_n502_), .A4(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n459_), .B1(new_n511_), .B2(new_n456_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n519_), .B(new_n522_), .Z(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n522_), .B(KEYINPUT15), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n519_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n519_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n530_), .A3(new_n524_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G113gat), .B(G141gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT76), .ZN(new_n534_));
  XOR2_X1   g333(.A(G169gat), .B(G197gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n532_), .B(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n512_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G85gat), .B(G92gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  INV_X1    g340(.A(G99gat), .ZN(new_n542_));
  INV_X1    g341(.A(G106gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT7), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT6), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(G99gat), .A3(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n541_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n550_), .B(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n545_), .B1(new_n554_), .B2(KEYINPUT67), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n550_), .B(KEYINPUT66), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n540_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n540_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n551_), .B1(new_n563_), .B2(KEYINPUT9), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(G85gat), .B2(G92gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT10), .B(G99gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT64), .ZN(new_n568_));
  OAI221_X1 g367(.A(new_n564_), .B1(new_n563_), .B2(new_n566_), .C1(new_n568_), .C2(G106gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n527_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n561_), .A2(new_n522_), .A3(new_n569_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(KEYINPUT70), .A3(new_n527_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n578_), .A2(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n573_), .A2(new_n581_), .A3(new_n586_), .A4(new_n582_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n592_), .B(KEYINPUT36), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n539_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n588_), .B2(KEYINPUT71), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n585_), .A2(new_n600_), .A3(new_n587_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n539_), .A3(new_n594_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n599_), .A2(new_n601_), .B1(new_n593_), .B2(new_n589_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(KEYINPUT72), .A3(new_n539_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n597_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n610_));
  XNOR2_X1  g409(.A(G57gat), .B(G64gat), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT11), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT11), .ZN(new_n613_));
  XOR2_X1   g412(.A(G71gat), .B(G78gat), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n613_), .A2(new_n614_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n570_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n561_), .A2(new_n617_), .A3(new_n569_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n610_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n570_), .A2(new_n618_), .B1(KEYINPUT68), .B2(KEYINPUT12), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n619_), .A2(new_n620_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT5), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n627_), .A2(new_n632_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n609_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n627_), .A2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n627_), .A2(new_n632_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT13), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(G127gat), .B(G155gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT16), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(KEYINPUT73), .A2(KEYINPUT17), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT17), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n519_), .B(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n617_), .ZN(new_n651_));
  MUX2_X1   g450(.A(new_n645_), .B(new_n648_), .S(new_n651_), .Z(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT74), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT74), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT75), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n608_), .A2(new_n639_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n538_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n446_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT38), .ZN(new_n662_));
  INV_X1    g461(.A(new_n459_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n502_), .A2(new_n510_), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n460_), .B(new_n407_), .C1(new_n495_), .C2(new_n498_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT102), .B1(new_n499_), .B2(new_n408_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n667_), .B2(new_n457_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n602_), .A2(new_n594_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n639_), .A2(new_n537_), .A3(new_n655_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n446_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n662_), .A3(new_n672_), .ZN(G1324gat));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  OAI21_X1  g473(.A(G8gat), .B1(new_n671_), .B2(new_n332_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n677_), .B(G8gat), .C1(new_n671_), .C2(new_n332_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(KEYINPUT39), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n538_), .A2(new_n515_), .A3(new_n331_), .A4(new_n658_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n676_), .B2(KEYINPUT39), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n674_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n684_), .A2(KEYINPUT40), .A3(new_n679_), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1325gat));
  OR3_X1    g485(.A1(new_n659_), .A2(G15gat), .A3(new_n456_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G15gat), .B1(new_n671_), .B2(new_n456_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n689_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1326gat));
  OR3_X1    g491(.A1(new_n659_), .A2(G22gat), .A3(new_n408_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G22gat), .B1(new_n671_), .B2(new_n408_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT42), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n597_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n607_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT72), .B1(new_n606_), .B2(new_n539_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n512_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n666_), .A2(new_n665_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n502_), .A2(new_n510_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n457_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n703_), .B(new_n608_), .C1(new_n706_), .C2(new_n459_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n702_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n537_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n638_), .A2(new_n635_), .A3(new_n657_), .A4(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT106), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n712_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n715_), .A2(KEYINPUT107), .A3(new_n490_), .A4(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G29gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT44), .B1(new_n708_), .B2(new_n712_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n714_), .B(new_n711_), .C1(new_n702_), .C2(new_n707_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n721_), .B2(new_n490_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n655_), .B(KEYINPUT75), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n669_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT108), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n639_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n538_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n446_), .A2(G29gat), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT109), .Z(new_n729_));
  OAI22_X1  g528(.A1(new_n718_), .A2(new_n722_), .B1(new_n727_), .B2(new_n729_), .ZN(G1328gat));
  NOR2_X1   g529(.A1(new_n332_), .A2(G36gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n727_), .A2(KEYINPUT45), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT45), .B1(new_n727_), .B2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n719_), .A2(new_n720_), .A3(new_n332_), .ZN(new_n736_));
  INV_X1    g535(.A(G36gat), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT46), .B(new_n735_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n715_), .A2(new_n331_), .A3(new_n716_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n739_), .A2(G36gat), .B1(new_n734_), .B2(new_n733_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n740_), .B2(new_n741_), .ZN(G1329gat));
  NOR2_X1   g541(.A1(new_n456_), .A2(new_n453_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n715_), .A2(new_n716_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n453_), .B1(new_n727_), .B2(new_n456_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(KEYINPUT47), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n745_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1330gat));
  INV_X1    g547(.A(new_n727_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G50gat), .B1(new_n749_), .B2(new_n407_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n407_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n721_), .B2(new_n751_), .ZN(G1331gat));
  NAND3_X1  g551(.A1(new_n701_), .A2(new_n639_), .A3(new_n723_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n512_), .A2(new_n709_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n490_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n668_), .A2(new_n669_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n639_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n709_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n723_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G57gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n490_), .B2(KEYINPUT112), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(KEYINPUT112), .B2(new_n765_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n759_), .B1(new_n764_), .B2(new_n767_), .ZN(G1332gat));
  INV_X1    g567(.A(G64gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n769_), .A3(new_n331_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n760_), .A2(new_n332_), .A3(new_n763_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G64gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G64gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT113), .B(new_n770_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n758_), .A2(new_n780_), .A3(new_n457_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n764_), .A2(new_n457_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G71gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  NOR2_X1   g585(.A1(new_n408_), .A2(G78gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n758_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n764_), .A2(new_n407_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G78gat), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n792_));
  AND2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n792_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n789_), .B1(new_n793_), .B2(new_n794_), .ZN(G1335gat));
  NAND2_X1  g594(.A1(new_n762_), .A2(new_n657_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n702_), .B2(new_n707_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798_), .B2(new_n446_), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n725_), .A2(new_n512_), .A3(new_n709_), .A4(new_n761_), .ZN(new_n800_));
  INV_X1    g599(.A(G85gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n490_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(G1336gat));
  OAI21_X1  g602(.A(G92gat), .B1(new_n798_), .B2(new_n332_), .ZN(new_n804_));
  INV_X1    g603(.A(G92gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n805_), .A3(new_n331_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1337gat));
  NOR2_X1   g606(.A1(new_n456_), .A2(new_n568_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n800_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n810_), .B(new_n542_), .C1(new_n797_), .C2(new_n457_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n796_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n708_), .A2(new_n457_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n813_), .B2(G99gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n809_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT51), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n809_), .C1(new_n811_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1338gat));
  NAND3_X1  g618(.A1(new_n800_), .A2(new_n543_), .A3(new_n407_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT52), .B(new_n543_), .C1(new_n797_), .C2(new_n407_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n708_), .A2(new_n407_), .A3(new_n812_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(G106gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT53), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n820_), .C1(new_n821_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n490_), .A2(new_n457_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n409_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT55), .B1(new_n625_), .B2(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(new_n610_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n626_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n622_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n623_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n623_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n835_), .A2(new_n842_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n631_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n523_), .A2(new_n524_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n528_), .A2(new_n530_), .A3(new_n525_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n536_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n532_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n536_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT119), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n845_), .A2(new_n856_), .A3(new_n631_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n834_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n847_), .A2(KEYINPUT58), .A3(new_n857_), .A4(new_n854_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n853_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n637_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n846_), .B2(KEYINPUT56), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n857_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n608_), .A2(new_n859_), .A3(new_n862_), .A4(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n853_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n637_), .A2(new_n709_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n856_), .A2(KEYINPUT118), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n846_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n845_), .A2(KEYINPUT118), .A3(new_n856_), .A4(new_n631_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n868_), .B1(new_n874_), .B2(new_n606_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n867_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n846_), .A2(new_n871_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n870_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n873_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n869_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT121), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n606_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(KEYINPUT57), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n723_), .B1(new_n876_), .B2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n701_), .A2(new_n537_), .A3(new_n761_), .A4(new_n723_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n833_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n874_), .A2(KEYINPUT121), .A3(new_n868_), .A4(new_n606_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n885_), .B1(new_n884_), .B2(KEYINPUT57), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n867_), .A2(new_n875_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n655_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n889_), .B(KEYINPUT54), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n832_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n892_), .B(new_n709_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G113gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n898_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n831_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n904_), .A2(G113gat), .A3(new_n537_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1340gat));
  OAI211_X1 g705(.A(new_n892_), .B(new_n639_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G120gat), .ZN(new_n908_));
  INV_X1    g707(.A(G120gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n761_), .B2(KEYINPUT60), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n909_), .B2(KEYINPUT60), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n899_), .B(new_n912_), .C1(new_n913_), .C2(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n908_), .A2(new_n914_), .ZN(G1341gat));
  AOI21_X1  g714(.A(G127gat), .B1(new_n899_), .B2(new_n723_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n657_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n898_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n904_), .A2(KEYINPUT59), .B1(new_n918_), .B2(new_n833_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT123), .B(G127gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n655_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n916_), .B1(new_n919_), .B2(new_n921_), .ZN(G1342gat));
  OAI211_X1 g721(.A(new_n892_), .B(new_n608_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G134gat), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n904_), .A2(G134gat), .A3(new_n669_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1343gat));
  NOR4_X1   g725(.A1(new_n331_), .A2(new_n408_), .A3(new_n446_), .A4(new_n457_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n903_), .A2(new_n709_), .A3(new_n927_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g728(.A1(new_n903_), .A2(new_n639_), .A3(new_n927_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g730(.A1(new_n903_), .A2(new_n723_), .A3(new_n927_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1346gat));
  NAND3_X1  g733(.A1(new_n903_), .A2(new_n608_), .A3(new_n927_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G162gat), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n669_), .A2(G162gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n903_), .A2(new_n927_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n332_), .A2(new_n458_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n709_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT124), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n408_), .B(new_n942_), .C1(new_n888_), .C2(new_n891_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n943_), .A2(new_n944_), .A3(G169gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n943_), .B2(G169gat), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n332_), .A2(new_n407_), .A3(new_n458_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n918_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n709_), .A2(new_n273_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT125), .Z(new_n950_));
  OAI22_X1  g749(.A1(new_n945_), .A2(new_n946_), .B1(new_n948_), .B2(new_n950_), .ZN(G1348gat));
  INV_X1    g750(.A(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n639_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n655_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n876_), .B2(new_n887_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n891_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(new_n407_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n639_), .A2(G176gat), .A3(new_n940_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n953_), .A2(new_n272_), .B1(new_n957_), .B2(new_n958_), .ZN(G1349gat));
  AOI21_X1  g758(.A(new_n655_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n903_), .A2(new_n408_), .A3(new_n723_), .A4(new_n940_), .ZN(new_n961_));
  AOI22_X1  g760(.A1(new_n952_), .A2(new_n960_), .B1(new_n961_), .B2(new_n236_), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n948_), .B2(new_n701_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n606_), .A2(new_n266_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n948_), .B2(new_n964_), .ZN(G1351gat));
  NOR3_X1   g764(.A1(new_n332_), .A2(new_n457_), .A3(new_n501_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n956_), .A2(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968_), .B2(new_n709_), .ZN(new_n969_));
  NOR4_X1   g768(.A1(new_n956_), .A2(new_n208_), .A3(new_n537_), .A4(new_n967_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1352gat));
  XNOR2_X1  g770(.A(KEYINPUT126), .B(G204gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n972_), .B1(new_n968_), .B2(new_n639_), .ZN(new_n973_));
  AND4_X1   g772(.A1(new_n639_), .A2(new_n903_), .A3(new_n966_), .A4(new_n972_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1353gat));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(KEYINPUT127), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n655_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n977_), .B1(new_n968_), .B2(new_n978_), .ZN(new_n979_));
  AND4_X1   g778(.A1(new_n903_), .A2(new_n966_), .A3(new_n978_), .A4(new_n977_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1354gat));
  NAND3_X1  g780(.A1(new_n968_), .A2(new_n224_), .A3(new_n606_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n956_), .A2(new_n701_), .A3(new_n967_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n982_), .B1(new_n224_), .B2(new_n983_), .ZN(G1355gat));
endmodule


