//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT79), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT24), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G190gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n213_), .A2(new_n215_), .A3(new_n217_), .A4(new_n219_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n210_), .A2(new_n211_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n211_), .B1(new_n210_), .B2(new_n220_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n207_), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT79), .B1(new_n204_), .B2(new_n205_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n221_), .A2(new_n222_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n212_), .A2(new_n216_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(KEYINPUT82), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(G169gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT22), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n205_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  AND4_X1   g042(.A1(new_n232_), .A2(new_n238_), .A3(new_n240_), .A4(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n203_), .B1(new_n230_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n222_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n210_), .A2(new_n220_), .A3(new_n211_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n226_), .A2(new_n228_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n232_), .A2(new_n238_), .A3(new_n240_), .A4(new_n243_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT83), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G43gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n252_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G15gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT85), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G113gat), .B(G120gat), .Z(new_n266_));
  OR3_X1    g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT31), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n261_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT88), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT1), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT87), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n283_), .A2(new_n280_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n269_), .B1(new_n300_), .B2(KEYINPUT93), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n284_), .A2(new_n289_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT93), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n304_), .A3(KEYINPUT4), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n300_), .A2(new_n308_), .A3(new_n269_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G29gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n301_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT33), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT95), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n310_), .A2(KEYINPUT33), .A3(new_n316_), .A4(new_n317_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n305_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n301_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n315_), .A3(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n327_), .A2(KEYINPUT90), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(KEYINPUT90), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT89), .B(G204gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(G197gat), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT21), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n328_), .A2(new_n329_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n333_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT21), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(KEYINPUT21), .A3(new_n338_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n328_), .A2(new_n329_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n336_), .A2(new_n340_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  INV_X1    g146(.A(new_n343_), .ZN(new_n348_));
  OAI22_X1  g147(.A1(new_n348_), .A2(new_n341_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n228_), .A2(new_n231_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT22), .B(G169gat), .Z(new_n351_));
  OAI211_X1 g150(.A(new_n350_), .B(new_n209_), .C1(G176gat), .C2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n223_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n353_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n220_), .A3(new_n210_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n349_), .B2(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n345_), .A2(new_n347_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n347_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n245_), .A2(new_n251_), .A3(new_n344_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n349_), .B2(new_n356_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n358_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n347_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n230_), .A2(new_n244_), .A3(new_n203_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(new_n249_), .B2(new_n250_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n349_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n357_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n359_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n368_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n318_), .A2(new_n380_), .A3(new_n319_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n321_), .A2(new_n326_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n310_), .A2(new_n317_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n315_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n318_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n372_), .A2(new_n377_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n360_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n359_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n385_), .B(new_n387_), .C1(new_n386_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n344_), .B1(KEYINPUT29), .B2(new_n300_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n302_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n302_), .B2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n398_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n398_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(KEYINPUT91), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n397_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n409_), .A2(KEYINPUT91), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n415_), .B(new_n396_), .C1(new_n409_), .C2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n393_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n385_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n370_), .B2(new_n378_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n369_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n372_), .A2(new_n368_), .A3(new_n377_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT27), .A3(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n417_), .A2(new_n420_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n274_), .B1(new_n419_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n347_), .B1(new_n345_), .B2(new_n357_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n368_), .B1(new_n428_), .B2(new_n388_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n370_), .A2(new_n429_), .A3(new_n421_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n369_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT27), .B1(new_n431_), .B2(new_n424_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT96), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n418_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT97), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT96), .B1(new_n430_), .B2(new_n432_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n422_), .A2(new_n434_), .A3(new_n425_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT97), .A3(new_n418_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n385_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n427_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT6), .ZN(new_n447_));
  OR3_X1    g246(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT65), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G85gat), .B(G92gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(KEYINPUT8), .A3(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(KEYINPUT9), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT10), .B(G99gat), .Z(new_n460_));
  INV_X1    g259(.A(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT64), .B(G85gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT9), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(G92gat), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n459_), .A2(new_n462_), .A3(new_n447_), .A4(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(new_n458_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT67), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT67), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n457_), .A2(new_n469_), .A3(new_n458_), .A4(new_n466_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n468_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G232gat), .A2(G233gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT34), .Z(new_n478_));
  INV_X1    g277(.A(KEYINPUT35), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n479_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT70), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n457_), .A2(new_n458_), .A3(new_n466_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n473_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n476_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n476_), .B2(new_n485_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G190gat), .B(G218gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G134gat), .B(G162gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT36), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(KEYINPUT36), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n488_), .B2(KEYINPUT71), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n476_), .A2(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n480_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n476_), .A2(new_n485_), .A3(new_n481_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(KEYINPUT71), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n494_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT99), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n488_), .A2(new_n492_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n488_), .A2(KEYINPUT71), .A3(new_n494_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n500_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT99), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n445_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT76), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G169gat), .B(G197gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n518_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G1gat), .B(G8gat), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n521_), .A2(new_n525_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n473_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT75), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT75), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n473_), .A3(new_n532_), .A4(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n475_), .A2(new_n529_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n517_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n473_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n516_), .B(new_n537_), .C1(new_n531_), .C2(new_n533_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n515_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT77), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n516_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n537_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n517_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n542_), .A2(new_n543_), .B1(new_n548_), .B2(new_n515_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n540_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT78), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(new_n515_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n468_), .A2(KEYINPUT12), .A3(new_n470_), .A4(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n566_), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(KEYINPUT66), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n467_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n484_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n484_), .A2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n569_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n575_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT13), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n556_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n529_), .B(new_n599_), .Z(new_n600_));
  AOI211_X1 g399(.A(new_n594_), .B(new_n598_), .C1(new_n600_), .C2(new_n564_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n564_), .B2(new_n600_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n600_), .A2(new_n573_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n598_), .B(KEYINPUT17), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n573_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n593_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT98), .Z(new_n610_));
  AND2_X1   g409(.A1(new_n511_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n202_), .B1(new_n611_), .B2(new_n385_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT100), .Z(new_n613_));
  INV_X1    g412(.A(KEYINPUT72), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n502_), .A2(new_n614_), .A3(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT72), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT72), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n508_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n608_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT74), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT97), .B1(new_n441_), .B2(new_n418_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n437_), .B(new_n417_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n444_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n274_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n417_), .B1(new_n382_), .B2(new_n392_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n426_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n593_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n624_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n202_), .A3(new_n385_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n613_), .A2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(new_n441_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n634_), .A2(new_n518_), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n511_), .A2(new_n638_), .A3(new_n610_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(G8gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n640_), .B2(G8gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n611_), .B2(new_n274_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n634_), .A2(new_n647_), .A3(new_n274_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n611_), .B2(new_n417_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n417_), .A2(new_n652_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT101), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n634_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(G1327gat));
  NAND2_X1  g457(.A1(new_n593_), .A2(new_n607_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n632_), .B2(new_n621_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT43), .B(new_n622_), .C1(new_n627_), .C2(new_n631_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT44), .B(new_n660_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(G29gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n420_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n445_), .B2(new_n622_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n632_), .A2(new_n661_), .A3(new_n621_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n659_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n670_));
  OAI211_X1 g469(.A(new_n664_), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n510_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n608_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n633_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n665_), .B1(new_n674_), .B2(new_n420_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(G1328gat));
  OAI211_X1 g475(.A(new_n664_), .B(new_n638_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n638_), .A2(KEYINPUT103), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n441_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n633_), .A2(new_n673_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n684_), .B(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n678_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n678_), .A2(KEYINPUT46), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  OAI21_X1  g491(.A(new_n664_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n274_), .A2(G43gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n674_), .A2(new_n628_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n693_), .A2(new_n694_), .B1(G43gat), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g496(.A1(new_n674_), .A2(G50gat), .A3(new_n418_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n664_), .B(new_n417_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT105), .B1(new_n699_), .B2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n592_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n555_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n445_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n624_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n385_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n705_), .A2(new_n607_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n511_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n420_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n682_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n511_), .A2(new_n715_), .A3(new_n710_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G64gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n707_), .A2(new_n723_), .A3(new_n274_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n711_), .A2(new_n628_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n723_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n711_), .B2(new_n418_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n707_), .A2(new_n733_), .A3(new_n417_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  AND2_X1   g534(.A1(new_n706_), .A2(new_n673_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n385_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n667_), .A2(new_n668_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n705_), .A2(new_n608_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT108), .Z(new_n741_));
  AND2_X1   g540(.A1(new_n385_), .A2(new_n463_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n737_), .B1(new_n741_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n736_), .B2(new_n638_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT109), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n715_), .A2(G92gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n741_), .B2(new_n746_), .ZN(G1337gat));
  NAND2_X1  g546(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n706_), .A2(new_n673_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n274_), .A2(new_n460_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n274_), .A3(new_n739_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(G99gat), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n736_), .A2(new_n461_), .A3(new_n417_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n417_), .B(new_n739_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G106gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n756_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  NAND3_X1  g564(.A1(new_n443_), .A2(new_n385_), .A3(new_n274_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n575_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n534_), .A2(new_n535_), .A3(new_n517_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n515_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n768_), .B(new_n769_), .C1(new_n517_), .C2(new_n546_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n539_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT113), .B1(new_n767_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n587_), .A2(new_n773_), .A3(new_n539_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n565_), .A2(new_n576_), .A3(new_n571_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n572_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n575_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n565_), .A2(new_n571_), .A3(new_n574_), .A4(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n585_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n775_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n775_), .B(KEYINPUT58), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n621_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n771_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n781_), .A2(new_n585_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT112), .A3(new_n791_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(new_n555_), .A3(new_n587_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n783_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n789_), .B1(new_n793_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n504_), .A2(new_n509_), .A3(KEYINPUT57), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n788_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n789_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n555_), .A3(new_n587_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT112), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n804_), .B2(new_n672_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n800_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n798_), .B2(new_n510_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(KEYINPUT57), .A3(new_n672_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .A4(new_n788_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n811_), .A3(new_n607_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n592_), .A2(new_n555_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(new_n615_), .A3(new_n608_), .A4(new_n620_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT54), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n766_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n555_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n766_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n766_), .A2(new_n818_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n814_), .B(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n808_), .A2(new_n810_), .A3(new_n788_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n607_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n608_), .B1(new_n825_), .B2(KEYINPUT114), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n828_), .B2(new_n811_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT115), .B(KEYINPUT59), .C1(new_n829_), .C2(new_n766_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n827_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n555_), .A2(new_n834_), .A3(G113gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n834_), .B2(G113gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n817_), .B1(new_n833_), .B2(new_n836_), .ZN(G1340gat));
  OAI21_X1  g636(.A(new_n592_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n816_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n703_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT60), .B2(new_n840_), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n839_), .A2(new_n840_), .B1(new_n841_), .B2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n816_), .B2(new_n608_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n608_), .A2(G127gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n833_), .B2(new_n846_), .ZN(G1342gat));
  AOI21_X1  g646(.A(G134gat), .B1(new_n816_), .B2(new_n510_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n621_), .A2(G134gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT118), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n833_), .B2(new_n850_), .ZN(G1343gat));
  NAND4_X1  g650(.A1(new_n682_), .A2(new_n385_), .A3(new_n417_), .A4(new_n628_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT119), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n555_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT120), .B(G141gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n592_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g658(.A1(new_n812_), .A2(new_n815_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n853_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n608_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT121), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n854_), .A2(new_n864_), .A3(new_n608_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(new_n854_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n870_), .A2(G162gat), .A3(new_n672_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G162gat), .B1(new_n870_), .B2(new_n622_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1347gat));
  AND3_X1   g672(.A1(new_n679_), .A2(new_n444_), .A3(new_n681_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n418_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n555_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n826_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n800_), .A2(new_n805_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n815_), .B1(new_n879_), .B2(new_n608_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n875_), .A2(new_n556_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n883_), .A3(G169gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n826_), .A2(new_n877_), .A3(new_n351_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT62), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n884_), .A2(new_n885_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n887_), .B(new_n888_), .C1(new_n890_), .C2(new_n891_), .ZN(G1348gat));
  NOR2_X1   g691(.A1(new_n829_), .A2(new_n417_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n874_), .A2(G176gat), .A3(new_n592_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n880_), .A2(new_n592_), .A3(new_n876_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n205_), .B2(new_n895_), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n880_), .A2(new_n876_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n607_), .B(new_n897_), .C1(new_n213_), .C2(new_n215_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n608_), .A3(new_n874_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n212_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n897_), .B2(new_n622_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n901_), .A2(KEYINPUT124), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(KEYINPUT124), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n510_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n902_), .A2(new_n903_), .B1(new_n897_), .B2(new_n904_), .ZN(G1351gat));
  NOR4_X1   g704(.A1(new_n682_), .A2(new_n385_), .A3(new_n418_), .A4(new_n274_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n860_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n332_), .B1(new_n907_), .B2(new_n556_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT126), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n910_), .B(new_n332_), .C1(new_n907_), .C2(new_n556_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n860_), .A2(G197gat), .A3(new_n555_), .A4(new_n906_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n913_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n909_), .A2(new_n911_), .B1(new_n914_), .B2(new_n915_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n907_), .A2(new_n703_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(G204gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n330_), .B2(new_n917_), .ZN(G1353gat));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920_));
  INV_X1    g719(.A(G211gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(new_n921_), .A3(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n860_), .A2(new_n608_), .A3(new_n906_), .A4(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT127), .B1(new_n920_), .B2(new_n921_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1354gat));
  OAI21_X1  g726(.A(G218gat), .B1(new_n907_), .B2(new_n622_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n672_), .A2(G218gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n907_), .B2(new_n929_), .ZN(G1355gat));
endmodule


