//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT23), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT79), .B(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT90), .Z(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT91), .Z(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n204_), .B1(KEYINPUT24), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n220_), .A2(KEYINPUT89), .B1(new_n213_), .B2(new_n214_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(KEYINPUT89), .B2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G204gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT84), .B1(new_n225_), .B2(G197gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(G197gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n225_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT21), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n227_), .B(KEYINPUT85), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(G197gat), .B2(new_n225_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n230_), .B(new_n231_), .C1(new_n233_), .C2(KEYINPUT21), .ZN(new_n234_));
  INV_X1    g033(.A(new_n231_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n224_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n213_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G169gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n206_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n205_), .A2(new_n209_), .A3(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G183gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT77), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n248_), .A3(G183gat), .ZN(new_n249_));
  INV_X1    g048(.A(G183gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT25), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n217_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n220_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n216_), .B1(new_n215_), .B2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n244_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n237_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT20), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT19), .ZN(new_n259_));
  NOR4_X1   g058(.A1(new_n239_), .A2(new_n256_), .A3(new_n257_), .A4(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n237_), .B2(new_n255_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n261_), .A2(KEYINPUT88), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(KEYINPUT88), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n224_), .A2(new_n238_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n265_), .B2(new_n259_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267_));
  INV_X1    g066(.A(G92gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT18), .B(G64gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(KEYINPUT27), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n265_), .A2(new_n259_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n259_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n256_), .A2(new_n257_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n237_), .A2(new_n223_), .A3(new_n211_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n271_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n265_), .A2(new_n259_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n271_), .B1(new_n281_), .B2(new_n260_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n284_));
  AOI22_X1  g083(.A1(new_n274_), .A2(new_n280_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT3), .Z(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT2), .Z(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n286_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n294_), .B2(new_n286_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n289_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n291_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n237_), .B1(KEYINPUT29), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G228gat), .A2(G233gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  XOR2_X1   g101(.A(G78gat), .B(G106gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n300_), .B(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT28), .ZN(new_n311_));
  XOR2_X1   g110(.A(G22gat), .B(G50gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT87), .A3(new_n307_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(KEYINPUT86), .A3(new_n307_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n285_), .A2(KEYINPUT96), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n283_), .A2(new_n284_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n273_), .A2(KEYINPUT27), .A3(new_n280_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT96), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n299_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n335_));
  AND3_X1   g134(.A1(new_n299_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n332_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(KEYINPUT92), .A3(KEYINPUT4), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n334_), .B1(new_n342_), .B2(new_n333_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  INV_X1    g143(.A(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G57gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n348_), .B(new_n334_), .C1(new_n342_), .C2(new_n333_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G71gat), .B(G99gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n255_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(new_n331_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT82), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT80), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n360_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n355_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n355_), .A2(new_n365_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n352_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n328_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n321_), .A2(new_n352_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n285_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n321_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n350_), .B(KEYINPUT33), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n342_), .A2(new_n333_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n333_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n349_), .B1(new_n337_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(KEYINPUT94), .A3(new_n377_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(new_n273_), .A3(new_n282_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n272_), .A2(KEYINPUT32), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n266_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n275_), .A2(new_n279_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n352_), .B(new_n385_), .C1(new_n386_), .C2(new_n384_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n373_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n368_), .B1(new_n372_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n370_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT15), .ZN(new_n391_));
  OR2_X1    g190(.A1(G29gat), .A2(G36gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G29gat), .A2(G36gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(G50gat), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G50gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(G29gat), .A2(G36gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G29gat), .A2(G36gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT69), .B(G43gat), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n394_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n391_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n394_), .A2(new_n398_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n399_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n394_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT15), .A3(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G99gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT10), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G99gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT64), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n345_), .A2(G92gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n268_), .A2(G85gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT9), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G99gat), .A2(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n345_), .A2(KEYINPUT9), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n268_), .A2(KEYINPUT65), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G92gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n419_), .A2(new_n422_), .A3(new_n427_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n425_), .A3(new_n426_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  XOR2_X1   g237(.A(G85gat), .B(G92gat), .Z(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n433_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n408_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n406_), .B2(new_n405_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G232gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n446_), .B(new_n451_), .C1(new_n444_), .C2(new_n443_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n450_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G190gat), .B(G218gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G134gat), .B(G162gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n459_), .B(KEYINPUT36), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n456_), .A2(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n467_), .B(new_n468_), .C1(new_n461_), .C2(new_n456_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G57gat), .A2(G64gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G57gat), .A2(G64gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT11), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G57gat), .ZN(new_n477_));
  INV_X1    g276(.A(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT11), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n473_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n471_), .B(KEYINPUT11), .C1(new_n475_), .C2(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G1gat), .A2(G8gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(G15gat), .A2(G22gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G15gat), .A2(G22gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(G1gat), .B2(G8gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n496_), .A2(new_n493_), .A3(new_n488_), .A4(new_n487_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n484_), .B(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n500_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT72), .B(KEYINPUT17), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G127gat), .B(G155gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G211gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT16), .B(G183gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n502_), .A2(new_n503_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT71), .B(KEYINPUT17), .Z(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n505_), .A2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n470_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n519_));
  INV_X1    g318(.A(new_n484_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n442_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n484_), .B(new_n433_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT12), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n442_), .A2(new_n524_), .A3(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT67), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  AOI211_X1 g329(.A(new_n529_), .B(new_n530_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n521_), .A2(new_n533_), .A3(new_n522_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n442_), .A2(KEYINPUT66), .A3(new_n520_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n225_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT5), .B(G176gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n519_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT13), .A3(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G169gat), .B(G197gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n402_), .A2(new_n407_), .A3(new_n498_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n495_), .B(new_n497_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT73), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n498_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(G229gat), .A3(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT74), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n562_), .B2(KEYINPUT75), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n551_), .A2(KEYINPUT75), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n561_), .B1(KEYINPUT74), .B2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n547_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n390_), .A2(new_n518_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n352_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(G1gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n202_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n569_), .B(KEYINPUT97), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(KEYINPUT98), .A3(new_n573_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(KEYINPUT38), .A3(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n390_), .A2(new_n568_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n462_), .A2(new_n465_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n517_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n572_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n575_), .A2(new_n577_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT99), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT99), .B1(new_n584_), .B2(new_n585_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n578_), .B(new_n583_), .C1(new_n587_), .C2(new_n588_), .ZN(G1324gat));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n285_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n486_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n576_), .A2(new_n486_), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n593_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1325gat));
  OAI21_X1  g401(.A(G15gat), .B1(new_n582_), .B2(new_n368_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT41), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT41), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n569_), .A2(G15gat), .A3(new_n368_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(G1326gat));
  OAI21_X1  g406(.A(G22gat), .B1(new_n582_), .B2(new_n321_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT42), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n321_), .A2(G22gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n569_), .B2(new_n610_), .ZN(G1327gat));
  INV_X1    g410(.A(new_n580_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n516_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n579_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(G29gat), .B1(new_n615_), .B2(new_n352_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n368_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n374_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n273_), .A2(new_n282_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n387_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n321_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n285_), .A2(new_n371_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n617_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n369_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n470_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n390_), .A2(new_n632_), .A3(KEYINPUT43), .A4(new_n470_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n631_), .A2(new_n633_), .A3(new_n517_), .A4(new_n568_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n636_), .A2(G29gat), .A3(new_n352_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n626_), .A2(new_n628_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n516_), .B1(new_n638_), .B2(new_n629_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n568_), .A4(new_n631_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n616_), .B1(new_n637_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n285_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(new_n640_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n285_), .A2(G36gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n615_), .A2(KEYINPUT45), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  INV_X1    g447(.A(new_n646_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n614_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n642_), .B1(new_n645_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT46), .ZN(G1329gat));
  XNOR2_X1  g452(.A(KEYINPUT104), .B(G43gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n636_), .A2(G43gat), .A3(new_n617_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n640_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n657_), .B(new_n659_), .ZN(G1330gat));
  AOI21_X1  g459(.A(G50gat), .B1(new_n615_), .B2(new_n373_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n395_), .B(new_n321_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(new_n640_), .ZN(G1331gat));
  AOI21_X1  g462(.A(new_n566_), .B1(new_n370_), .B2(new_n389_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n547_), .A3(new_n581_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(new_n477_), .A3(new_n572_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n547_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n390_), .A2(new_n567_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n518_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT107), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n352_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n666_), .B1(new_n675_), .B2(new_n477_), .ZN(G1332gat));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n478_), .A3(new_n591_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G64gat), .B1(new_n665_), .B2(new_n285_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n681_), .A3(new_n617_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G71gat), .B1(new_n665_), .B2(new_n368_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT49), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1334gat));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n674_), .A2(new_n686_), .A3(new_n373_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G78gat), .B1(new_n665_), .B2(new_n321_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT50), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1335gat));
  NOR2_X1   g489(.A1(new_n667_), .A2(new_n566_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n631_), .A2(new_n633_), .A3(new_n517_), .A4(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n345_), .A3(new_n572_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n672_), .A2(new_n613_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n352_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n345_), .ZN(G1336gat));
  AOI21_X1  g495(.A(G92gat), .B1(new_n694_), .B2(new_n591_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n692_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n591_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(G1337gat));
  AOI21_X1  g499(.A(new_n368_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n670_), .A2(new_n613_), .A3(new_n671_), .A4(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT108), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n617_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n704_), .A2(G99gat), .B1(new_n705_), .B2(KEYINPUT51), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT51), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n703_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1338gat));
  NAND4_X1  g510(.A1(new_n672_), .A2(new_n418_), .A3(new_n373_), .A4(new_n613_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n698_), .A2(new_n373_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G106gat), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n713_), .B(G106gat), .C1(new_n692_), .C2(new_n321_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n712_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT53), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT53), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n712_), .B(new_n720_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1339gat));
  XOR2_X1   g521(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n527_), .A2(KEYINPUT111), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n523_), .A2(new_n525_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n527_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n532_), .B2(new_n727_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n724_), .B1(new_n732_), .B2(new_n540_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n522_), .A2(KEYINPUT12), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n437_), .A2(new_n439_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT8), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n484_), .B1(new_n738_), .B2(new_n433_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n734_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n525_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n527_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n529_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n526_), .A2(KEYINPUT67), .A3(new_n527_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n727_), .A3(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n729_), .A2(new_n730_), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n724_), .B(new_n540_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n733_), .B1(new_n747_), .B2(KEYINPUT116), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n540_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n749_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n557_), .A2(new_n560_), .A3(new_n550_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n555_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT113), .B1(new_n753_), .B2(new_n550_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n753_), .A2(KEYINPUT113), .A3(new_n550_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n752_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .A3(new_n541_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n760_), .A2(new_n761_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n542_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n723_), .B1(new_n751_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n466_), .A2(new_n469_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n748_), .A2(new_n750_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n470_), .B(new_n771_), .C1(new_n772_), .C2(new_n723_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n751_), .A2(KEYINPUT58), .A3(new_n767_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n770_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n765_), .B1(new_n545_), .B2(new_n541_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n747_), .A3(KEYINPUT112), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n566_), .B(new_n541_), .C1(new_n733_), .C2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n566_), .A2(new_n541_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n779_), .B2(KEYINPUT112), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n733_), .A2(new_n788_), .A3(new_n781_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n777_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n790_), .B2(new_n580_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n784_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n516_), .B1(new_n776_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n566_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n544_), .A2(new_n546_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n769_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n797_), .B2(new_n769_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n793_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n769_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT54), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n799_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n784_), .A2(new_n791_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n470_), .B1(new_n772_), .B2(new_n723_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n774_), .B1(new_n809_), .B2(KEYINPUT118), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(new_n773_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n806_), .B(new_n807_), .C1(new_n811_), .C2(new_n516_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n803_), .A2(new_n812_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n572_), .B(new_n368_), .C1(new_n322_), .C2(new_n327_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n566_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n806_), .B1(new_n811_), .B2(new_n516_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n814_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n815_), .B2(KEYINPUT59), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n566_), .A2(G113gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n667_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n816_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n824_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n821_), .A2(new_n547_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n824_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n816_), .B2(new_n516_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n516_), .A2(G127gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n821_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n816_), .B2(new_n580_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n470_), .A2(G134gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT121), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n821_), .B2(new_n834_), .ZN(G1343gat));
  NOR3_X1   g634(.A1(new_n591_), .A2(new_n572_), .A3(new_n321_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n813_), .A2(new_n368_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n566_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n547_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g641(.A1(new_n837_), .A2(new_n517_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1346gat));
  INV_X1    g644(.A(G162gat), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n837_), .A2(new_n846_), .A3(new_n769_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n838_), .A2(new_n580_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1347gat));
  NOR3_X1   g648(.A1(new_n285_), .A2(new_n373_), .A3(new_n624_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n818_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G169gat), .B1(new_n852_), .B2(new_n567_), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n853_), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n853_), .B2(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(KEYINPUT62), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n566_), .A3(new_n207_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1348gat));
  AND2_X1   g658(.A1(new_n813_), .A2(new_n850_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n667_), .A2(new_n214_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n851_), .A2(new_n547_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n860_), .A2(new_n861_), .B1(new_n206_), .B2(new_n862_), .ZN(G1349gat));
  AOI21_X1  g662(.A(G183gat), .B1(new_n860_), .B2(new_n516_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n517_), .A2(new_n218_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n851_), .B2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n852_), .B2(new_n769_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n851_), .A2(new_n580_), .A3(new_n217_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1351gat));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n591_), .A2(new_n371_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n803_), .A2(new_n368_), .A3(new_n812_), .A4(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n567_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n870_), .B1(new_n874_), .B2(G197gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  INV_X1    g675(.A(G197gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n876_), .A2(KEYINPUT123), .A3(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n875_), .B(new_n878_), .C1(new_n876_), .C2(new_n877_), .ZN(G1352gat));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n873_), .A2(new_n667_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n225_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n873_), .B2(new_n667_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G204gat), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n873_), .A2(new_n883_), .A3(new_n667_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n889_), .A2(new_n880_), .A3(G204gat), .A4(new_n884_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n887_), .A2(new_n888_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n888_), .B1(new_n887_), .B2(new_n890_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1353gat));
  XNOR2_X1  g692(.A(KEYINPUT63), .B(G211gat), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n873_), .A2(new_n517_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT127), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n895_), .A2(KEYINPUT127), .ZN(new_n897_));
  INV_X1    g696(.A(new_n873_), .ZN(new_n898_));
  AOI211_X1 g697(.A(KEYINPUT63), .B(G211gat), .C1(new_n898_), .C2(new_n516_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n897_), .B2(new_n899_), .ZN(G1354gat));
  INV_X1    g699(.A(G218gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n873_), .A2(new_n901_), .A3(new_n769_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n580_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n901_), .B2(new_n903_), .ZN(G1355gat));
endmodule


