//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT21), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n203_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n204_), .A2(new_n208_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n202_), .B1(new_n211_), .B2(new_n206_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214_));
  AND2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(KEYINPUT86), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n220_), .B(new_n221_), .C1(new_n222_), .C2(KEYINPUT2), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n217_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n217_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n214_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(G228gat), .B(G233gat), .C1(new_n213_), .C2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n231_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT87), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n227_), .A2(new_n236_), .A3(new_n231_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n214_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n210_), .A2(new_n212_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n233_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n237_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT29), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(new_n241_), .A3(new_n243_), .A4(new_n240_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n246_), .B1(new_n252_), .B2(new_n233_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT91), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n247_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n246_), .A3(new_n233_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n235_), .A2(new_n214_), .A3(new_n237_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G22gat), .B(G50gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n260_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n262_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n258_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n270_), .A2(new_n256_), .A3(new_n257_), .A4(new_n255_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT19), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G176gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT23), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n276_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(KEYINPUT92), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(KEYINPUT92), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(KEYINPUT82), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n280_), .A2(new_n292_), .A3(KEYINPUT23), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n285_), .A2(KEYINPUT24), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G190gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .A4(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n213_), .A2(new_n284_), .A3(new_n298_), .ZN(new_n299_));
  OAI221_X1 g098(.A(new_n293_), .B1(G183gat), .B2(G190gat), .C1(new_n281_), .C2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n279_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n302_));
  INV_X1    g101(.A(G190gat), .ZN(new_n303_));
  OR3_X1    g102(.A1(new_n303_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT26), .B1(new_n303_), .B2(KEYINPUT81), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n295_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n281_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n243_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n274_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n298_), .A2(new_n284_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n243_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n274_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n213_), .A2(new_n301_), .A3(new_n307_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n315_), .A2(new_n317_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n274_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n324_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n299_), .A2(new_n309_), .A3(KEYINPUT20), .A4(new_n316_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(KEYINPUT27), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n272_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT98), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT85), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n344_), .A2(new_n345_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n249_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n346_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n227_), .A2(new_n351_), .A3(new_n231_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n343_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT4), .B1(new_n249_), .B2(new_n349_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n342_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n341_), .A3(new_n352_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n355_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G15gat), .B(G43gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT83), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n367_), .B(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n308_), .B(KEYINPUT30), .Z(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(KEYINPUT84), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(KEYINPUT84), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  XOR2_X1   g173(.A(new_n349_), .B(KEYINPUT31), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n272_), .A2(KEYINPUT98), .A3(new_n337_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n340_), .A2(new_n364_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT99), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT98), .B1(new_n272_), .B2(new_n337_), .ZN(new_n382_));
  AOI211_X1 g181(.A(new_n339_), .B(new_n336_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n384_), .A2(KEYINPUT99), .A3(new_n364_), .A4(new_n377_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n328_), .A2(KEYINPUT32), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n319_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT96), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n327_), .A2(new_n329_), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n362_), .A2(new_n363_), .B1(new_n390_), .B2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n355_), .A2(new_n356_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n333_), .A2(new_n334_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n355_), .A2(KEYINPUT33), .A3(new_n356_), .A4(new_n361_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n341_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n353_), .A2(new_n354_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n341_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n361_), .B1(new_n400_), .B2(KEYINPUT33), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n389_), .A2(new_n391_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n272_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT97), .ZN(new_n404_));
  INV_X1    g203(.A(new_n272_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n364_), .A3(new_n337_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n402_), .A2(new_n407_), .A3(new_n272_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n376_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n386_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT12), .ZN(new_n412_));
  XOR2_X1   g211(.A(G85gat), .B(G92gat), .Z(new_n413_));
  OR2_X1    g212(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n414_));
  NAND2_X1  g213(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G99gat), .A2(G106gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT6), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n414_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT10), .B(G99gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(G106gat), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n416_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n424_));
  NOR4_X1   g223(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT66), .A2(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n424_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT66), .ZN(new_n431_));
  INV_X1    g230(.A(G99gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT7), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT68), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n436_), .A3(new_n418_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n413_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT69), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n440_), .A3(new_n413_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(KEYINPUT8), .A3(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n425_), .A2(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n418_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT8), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n447_), .A3(new_n418_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n413_), .A4(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n423_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G64gat), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n453_));
  XOR2_X1   g252(.A(G71gat), .B(G78gat), .Z(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n453_), .A2(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n412_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n423_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n437_), .A2(new_n440_), .A3(new_n413_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n440_), .B1(new_n437_), .B2(new_n413_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n446_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n449_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n457_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT12), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G230gat), .A2(G233gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT64), .Z(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT71), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n458_), .A2(new_n466_), .A3(new_n469_), .A4(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n450_), .A2(new_n457_), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n465_), .B(new_n423_), .C1(new_n442_), .C2(new_n449_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n468_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT70), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n479_), .B(new_n468_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G176gat), .B(G204gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G120gat), .B(G148gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n474_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n490_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n487_), .B1(new_n474_), .B2(new_n481_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT74), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT74), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT77), .B(G8gat), .Z(new_n502_));
  AND2_X1   g301(.A1(new_n502_), .A2(KEYINPUT14), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G1gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n503_), .A2(new_n505_), .B1(new_n507_), .B2(G1gat), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(G8gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(G8gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT78), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n457_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n512_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G127gat), .B(G155gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n521_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G232gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT34), .ZN(new_n534_));
  XOR2_X1   g333(.A(G43gat), .B(G50gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT15), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n450_), .A2(new_n538_), .ZN(new_n539_));
  AOI211_X1 g338(.A(new_n423_), .B(new_n537_), .C1(new_n442_), .C2(new_n449_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT35), .B(new_n534_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n464_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n537_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n450_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n534_), .A2(KEYINPUT35), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n534_), .A2(KEYINPUT35), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_));
  AOI211_X1 g347(.A(new_n530_), .B(new_n532_), .C1(new_n541_), .C2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n529_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT76), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n541_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT37), .B1(new_n549_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n541_), .A2(new_n548_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n530_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n531_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n553_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n526_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n511_), .A2(new_n538_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n511_), .B2(new_n544_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n511_), .B(new_n544_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT80), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AND4_X1   g377(.A1(new_n411_), .A2(new_n501_), .A3(new_n561_), .A4(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G1gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n364_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n501_), .A2(new_n576_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n558_), .A2(new_n553_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n586_), .A2(new_n526_), .A3(new_n588_), .A4(new_n411_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n364_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(G1324gat));
  NAND3_X1  g390(.A1(new_n579_), .A2(new_n502_), .A3(new_n336_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G8gat), .B1(new_n589_), .B2(new_n337_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(G1325gat));
  OAI21_X1  g397(.A(G15gat), .B1(new_n589_), .B2(new_n376_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT41), .Z(new_n600_));
  INV_X1    g399(.A(G15gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n579_), .A2(new_n601_), .A3(new_n377_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(G1326gat));
  INV_X1    g402(.A(G22gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n272_), .B(KEYINPUT101), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n579_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G22gat), .B1(new_n589_), .B2(new_n605_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1327gat));
  NOR2_X1   g412(.A1(new_n526_), .A2(new_n588_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n411_), .A2(new_n501_), .A3(new_n578_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n616_), .B2(new_n581_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n526_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n555_), .A2(new_n560_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n411_), .B2(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n381_), .A2(new_n385_), .B1(new_n376_), .B2(new_n409_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(KEYINPUT43), .A3(new_n620_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n618_), .B(new_n586_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n627_), .A2(G29gat), .A3(new_n581_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n411_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT43), .B1(new_n623_), .B2(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n631_), .A2(KEYINPUT44), .A3(new_n618_), .A4(new_n586_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n617_), .B1(new_n628_), .B2(new_n632_), .ZN(G1328gat));
  XNOR2_X1  g432(.A(new_n336_), .B(KEYINPUT103), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n615_), .A2(G36gat), .A3(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n637_));
  XOR2_X1   g436(.A(new_n636_), .B(new_n637_), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n336_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n585_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT44), .B1(new_n640_), .B2(new_n618_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G36gat), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n642_), .A3(KEYINPUT46), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  INV_X1    g446(.A(KEYINPUT47), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  INV_X1    g448(.A(G43gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n650_), .B1(new_n615_), .B2(new_n376_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n376_), .A2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n632_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n649_), .B(new_n651_), .C1(new_n653_), .C2(new_n641_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n627_), .A2(new_n632_), .A3(new_n652_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n656_), .B2(new_n651_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n648_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n653_), .B2(new_n641_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(KEYINPUT47), .A3(new_n654_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n616_), .B2(new_n606_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n627_), .A2(G50gat), .A3(new_n632_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n405_), .ZN(G1331gat));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(new_n576_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n411_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT106), .B1(new_n623_), .B2(new_n576_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n501_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n561_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n364_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(KEYINPUT107), .A3(new_n561_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G57gat), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n677_), .B(G57gat), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n501_), .A2(new_n618_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n679_), .A2(new_n411_), .A3(new_n588_), .A4(new_n577_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n680_), .A2(KEYINPUT109), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(KEYINPUT109), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n681_), .A2(G57gat), .A3(new_n581_), .A4(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n676_), .A2(new_n678_), .A3(new_n685_), .ZN(G1332gat));
  OR3_X1    g485(.A1(new_n671_), .A2(G64gat), .A3(new_n635_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n681_), .A2(new_n634_), .A3(new_n682_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G64gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G64gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1333gat));
  OR3_X1    g491(.A1(new_n671_), .A2(G71gat), .A3(new_n376_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n681_), .A2(new_n377_), .A3(new_n682_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G71gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1334gat));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n606_), .A3(new_n682_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(G78gat), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G78gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n605_), .A2(G78gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT112), .Z(new_n704_));
  OAI22_X1  g503(.A1(new_n701_), .A2(new_n702_), .B1(new_n671_), .B2(new_n704_), .ZN(G1335gat));
  AND2_X1   g504(.A1(new_n670_), .A2(new_n614_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n581_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n501_), .A2(new_n526_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n631_), .A2(new_n667_), .A3(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT113), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT113), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n364_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n712_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n706_), .B2(new_n336_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n635_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n718_));
  INV_X1    g517(.A(new_n421_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n706_), .A2(new_n719_), .A3(new_n377_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G99gat), .B1(new_n709_), .B2(new_n376_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT115), .Z(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n722_), .B(new_n725_), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n428_), .A3(new_n405_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n631_), .A2(new_n708_), .A3(new_n405_), .A4(new_n667_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G106gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G106gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(G113gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT59), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(KEYINPUT118), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n494_), .A2(new_n495_), .A3(new_n491_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n497_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n561_), .B(new_n577_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT116), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n498_), .A2(new_n742_), .A3(new_n561_), .A4(new_n577_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n741_), .A2(new_n743_), .A3(KEYINPUT54), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT54), .B1(new_n741_), .B2(new_n743_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n490_), .A2(new_n576_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT55), .B1(new_n471_), .B2(new_n473_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n466_), .A2(new_n458_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n468_), .B1(new_n749_), .B2(new_n476_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n458_), .A2(new_n466_), .A3(new_n469_), .A4(KEYINPUT55), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n488_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT56), .B(new_n488_), .C1(new_n748_), .C2(new_n752_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n747_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n563_), .A2(new_n567_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n566_), .A2(new_n564_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n572_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n575_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n588_), .B1(new_n757_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT57), .B(new_n588_), .C1(new_n757_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n490_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT117), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n490_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n755_), .A2(new_n756_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(KEYINPUT58), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT58), .B1(new_n773_), .B2(new_n774_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n620_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n618_), .B1(new_n767_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n364_), .B1(new_n746_), .B2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n382_), .A2(new_n383_), .A3(new_n376_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n737_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n746_), .A2(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n581_), .A3(new_n780_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n735_), .A2(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n781_), .B1(new_n785_), .B2(new_n737_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n734_), .B1(new_n786_), .B2(new_n578_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n783_), .A2(G113gat), .A3(new_n667_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT119), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n736_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n779_), .A2(new_n780_), .B1(KEYINPUT118), .B2(new_n735_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n736_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n577_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  INV_X1    g593(.A(new_n788_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n789_), .A2(new_n796_), .ZN(G1340gat));
  OAI21_X1  g596(.A(KEYINPUT120), .B1(new_n792_), .B2(new_n501_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  INV_X1    g598(.A(new_n501_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n801_), .A3(G120gat), .ZN(new_n802_));
  INV_X1    g601(.A(new_n783_), .ZN(new_n803_));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n501_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n803_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n804_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(G1341gat));
  AOI21_X1  g606(.A(G127gat), .B1(new_n803_), .B2(new_n526_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n526_), .A2(G127gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n786_), .B2(new_n809_), .ZN(G1342gat));
  AOI21_X1  g609(.A(G134gat), .B1(new_n803_), .B2(new_n587_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT121), .B(G134gat), .Z(new_n812_));
  NOR2_X1   g611(.A1(new_n620_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n786_), .B2(new_n813_), .ZN(G1343gat));
  AND2_X1   g613(.A1(new_n779_), .A2(new_n635_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n377_), .A2(new_n272_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n667_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT122), .B(G141gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1344gat));
  INV_X1    g619(.A(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n800_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g622(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n817_), .B2(new_n618_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n815_), .A2(new_n526_), .A3(new_n816_), .A4(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n829_), .A3(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1346gat));
  AND3_X1   g632(.A1(new_n821_), .A2(G162gat), .A3(new_n621_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G162gat), .B1(new_n821_), .B2(new_n587_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1347gat));
  AOI21_X1  g635(.A(new_n606_), .B1(new_n746_), .B2(new_n778_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n635_), .A2(new_n581_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n377_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT125), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n667_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n278_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n275_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT62), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(KEYINPUT62), .B2(new_n845_), .ZN(G1348gat));
  INV_X1    g646(.A(new_n842_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G176gat), .B1(new_n848_), .B2(new_n800_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n405_), .B1(new_n746_), .B2(new_n778_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n840_), .A2(new_n276_), .A3(new_n501_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n840_), .A2(new_n618_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G183gat), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n840_), .A2(new_n618_), .A3(new_n295_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n837_), .B2(new_n855_), .ZN(G1350gat));
  NAND3_X1  g655(.A1(new_n848_), .A2(new_n587_), .A3(new_n296_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n621_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n858_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT126), .B1(new_n858_), .B2(G190gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(G1351gat));
  AND2_X1   g660(.A1(new_n782_), .A2(new_n816_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n838_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n576_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n800_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g667(.A1(new_n863_), .A2(new_n618_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  AND2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n869_), .B2(new_n870_), .ZN(G1354gat));
  OR3_X1    g672(.A1(new_n863_), .A2(KEYINPUT127), .A3(new_n588_), .ZN(new_n874_));
  INV_X1    g673(.A(G218gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT127), .B1(new_n863_), .B2(new_n588_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n864_), .A2(G218gat), .A3(new_n621_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1355gat));
endmodule


