//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT73), .Z(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT8), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n215_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT66), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(new_n215_), .C1(new_n220_), .C2(new_n226_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n213_), .A2(new_n214_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n217_), .A2(new_n219_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n226_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT67), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n228_), .B(new_n230_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G29gat), .B(G36gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G43gat), .B(G50gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n223_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n220_), .B1(KEYINPUT64), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n214_), .B1(new_n213_), .B2(KEYINPUT9), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n247_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n246_), .B(new_n251_), .C1(KEYINPUT64), .C2(new_n245_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n239_), .A2(new_n242_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n228_), .A2(new_n230_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n234_), .A2(new_n233_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n224_), .A2(new_n225_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n236_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n238_), .B1(new_n259_), .B2(new_n231_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n242_), .B(KEYINPUT15), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT74), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n265_), .A3(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT75), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n255_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(KEYINPUT75), .A3(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n211_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n267_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n255_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n211_), .ZN(new_n274_));
  OAI22_X1  g073(.A1(new_n271_), .A2(KEYINPUT76), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276_));
  AOI211_X1 g075(.A(new_n276_), .B(new_n211_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n206_), .B(new_n207_), .C1(new_n275_), .C2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n272_), .A2(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n268_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n211_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n279_), .B1(new_n283_), .B2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(KEYINPUT76), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n205_), .A3(new_n204_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n278_), .B2(new_n286_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G183gat), .B(G211gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT80), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT17), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT70), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT78), .ZN(new_n305_));
  XOR2_X1   g104(.A(G15gat), .B(G22gat), .Z(new_n306_));
  NAND2_X1  g105(.A1(G1gat), .A2(G8gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(KEYINPUT14), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n305_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G64gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G78gat), .Z(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n314_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n311_), .B(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n303_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n299_), .A2(new_n302_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n293_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT81), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n261_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n261_), .A2(KEYINPUT70), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT12), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n261_), .B(new_n327_), .C1(KEYINPUT70), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n319_), .B(new_n252_), .C1(new_n256_), .C2(new_n260_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT71), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n338_), .A3(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n239_), .A2(KEYINPUT68), .A3(new_n319_), .A4(new_n252_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n328_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n346_));
  INV_X1    g145(.A(new_n335_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n341_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G120gat), .B(G148gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT5), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G176gat), .B(G204gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n341_), .B(new_n356_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT13), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(KEYINPUT13), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT72), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT87), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT2), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(KEYINPUT85), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(KEYINPUT85), .B2(new_n382_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n377_), .A2(new_n385_), .A3(KEYINPUT1), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n377_), .B1(new_n378_), .B2(KEYINPUT1), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n377_), .B2(KEYINPUT1), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n384_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n380_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G127gat), .B(G134gat), .Z(new_n392_));
  XOR2_X1   g191(.A(G113gat), .B(G120gat), .Z(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n380_), .A3(new_n390_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(KEYINPUT4), .A3(new_n397_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n391_), .A2(new_n403_), .A3(new_n394_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n368_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT101), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT18), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT19), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT82), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT24), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT26), .B(G190gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT25), .B(G183gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(KEYINPUT23), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G169gat), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n417_), .A2(KEYINPUT24), .A3(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n418_), .A2(new_n421_), .A3(new_n426_), .A4(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT84), .B1(new_n427_), .B2(KEYINPUT22), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n428_), .B(new_n433_), .C1(new_n434_), .C2(KEYINPUT84), .ZN(new_n435_));
  INV_X1    g234(.A(new_n422_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n424_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(KEYINPUT23), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n430_), .B(new_n435_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n432_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G211gat), .B(G218gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT92), .B(G197gat), .ZN(new_n444_));
  INV_X1    g243(.A(G204gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT21), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(G197gat), .B2(G204gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n443_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(G197gat), .A2(G204gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n444_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(G204gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n449_), .B1(new_n452_), .B2(KEYINPUT21), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(KEYINPUT21), .A3(new_n443_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT93), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(KEYINPUT93), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n442_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n439_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT24), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n416_), .A2(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n459_), .A2(new_n431_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n420_), .B(KEYINPUT97), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n419_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n425_), .A2(new_n440_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n429_), .B1(new_n434_), .B2(new_n428_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n462_), .A2(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n453_), .A2(new_n454_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n415_), .B1(new_n458_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT98), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n472_), .B(new_n415_), .C1(new_n458_), .C2(new_n469_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n456_), .A2(new_n457_), .A3(new_n442_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n415_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT20), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n413_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n413_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n477_), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n479_), .B(new_n480_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT33), .B(new_n368_), .C1(new_n401_), .C2(new_n405_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT99), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n398_), .A2(new_n400_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n402_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n368_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n409_), .A2(new_n482_), .A3(new_n484_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n477_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n465_), .A2(new_n466_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n463_), .A2(new_n419_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n459_), .A2(new_n431_), .A3(new_n461_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT102), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n468_), .A2(KEYINPUT95), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n455_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n492_), .B(KEYINPUT102), .C1(new_n493_), .C2(new_n494_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n475_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT103), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n415_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n503_), .B2(new_n415_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n458_), .A2(new_n469_), .A3(new_n415_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n491_), .B1(new_n508_), .B2(new_n490_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n401_), .A2(new_n405_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n487_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT104), .A3(new_n406_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT104), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(new_n487_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT105), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n512_), .A2(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n490_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n506_), .A2(new_n507_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n505_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT105), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n520_), .A3(new_n521_), .A4(new_n491_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n489_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G228gat), .A2(G233gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n456_), .A2(new_n457_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n391_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n529_));
  AND4_X1   g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(KEYINPUT94), .A2(new_n526_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n526_), .A2(KEYINPUT94), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n524_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT96), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G22gat), .B(G50gat), .Z(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT28), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n391_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n539_), .A2(KEYINPUT90), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n391_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n538_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT90), .B1(new_n539_), .B2(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n537_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n542_), .A3(new_n538_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT96), .B1(new_n530_), .B2(new_n533_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G78gat), .B(G106gat), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n536_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n554_), .A3(new_n535_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n517_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n482_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n564_));
  OAI21_X1  g363(.A(new_n479_), .B1(new_n519_), .B2(new_n505_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT27), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n481_), .A2(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n563_), .A2(new_n564_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n523_), .A2(new_n561_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G71gat), .B(G99gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G43gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n442_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n396_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G227gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(G15gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT30), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT31), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n573_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n561_), .A2(new_n568_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n515_), .A2(new_n579_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n569_), .A2(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n309_), .B(new_n242_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT15), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n242_), .B(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(new_n309_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n309_), .A2(new_n242_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G169gat), .B(G197gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n582_), .A2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n326_), .A2(new_n364_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(G1gat), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n517_), .A2(KEYINPUT107), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n517_), .A2(KEYINPUT107), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n582_), .A2(new_n287_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n362_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n599_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n324_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n515_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n606_), .A2(new_n607_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n616_), .A3(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(G8gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n568_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n601_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n620_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n623_), .B2(G8gat), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT39), .B(new_n619_), .C1(new_n614_), .C2(new_n620_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(new_n579_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G15gat), .B1(new_n615_), .B2(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n601_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n561_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n614_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n601_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1327gat));
  AND2_X1   g440(.A1(new_n278_), .A2(new_n286_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n612_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT109), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n362_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n600_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n517_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n611_), .A2(new_n324_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(new_n293_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n582_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n582_), .B2(new_n650_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n605_), .A2(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n647_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n620_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n568_), .A2(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n600_), .A2(new_n645_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n661_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT46), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n660_), .B2(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(KEYINPUT110), .A3(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n669_), .A2(new_n672_), .ZN(G1329gat));
  NAND3_X1  g472(.A1(new_n657_), .A2(G43gat), .A3(new_n579_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n646_), .A2(new_n579_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(G43gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT47), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1330gat));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n646_), .A2(new_n682_), .A3(new_n636_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n657_), .A2(KEYINPUT111), .A3(new_n636_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G50gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT111), .B1(new_n657_), .B2(new_n636_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n612_), .A2(new_n599_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n363_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n609_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G57gat), .B1(new_n691_), .B2(new_n515_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n599_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n582_), .A2(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n326_), .A2(new_n362_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G57gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n605_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n692_), .A2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(G64gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n690_), .B2(new_n620_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n699_), .A3(new_n620_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1333gat));
  INV_X1    g503(.A(G71gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n690_), .B2(new_n579_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n705_), .A3(new_n579_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1334gat));
  INV_X1    g509(.A(G78gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n690_), .B2(new_n636_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT50), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n695_), .A2(new_n711_), .A3(new_n636_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n644_), .A2(new_n364_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n694_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G85gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n605_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n651_), .A2(new_n652_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n610_), .A2(new_n324_), .A3(new_n599_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n517_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n724_), .B2(new_n719_), .ZN(G1336gat));
  INV_X1    g524(.A(G92gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n726_), .A3(new_n620_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n723_), .A2(new_n620_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n726_), .ZN(G1337gat));
  AOI21_X1  g528(.A(new_n222_), .B1(new_n723_), .B2(new_n579_), .ZN(new_n730_));
  AND4_X1   g529(.A1(new_n243_), .A2(new_n718_), .A3(new_n244_), .A4(new_n579_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n730_), .A2(KEYINPUT51), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT51), .B1(new_n730_), .B2(new_n731_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n223_), .A3(new_n636_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n721_), .A2(new_n636_), .A3(new_n722_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n223_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n735_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT119), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n332_), .A2(new_n330_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n343_), .A2(new_n344_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n747_), .A2(KEYINPUT55), .B1(new_n749_), .B2(new_n335_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n333_), .A2(new_n340_), .A3(KEYINPUT55), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n354_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT56), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n354_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n583_), .A2(new_n584_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n589_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n596_), .A3(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n357_), .A2(new_n598_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n755_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n753_), .A2(new_n759_), .A3(KEYINPUT58), .A4(new_n755_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n287_), .A2(new_n288_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n291_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n357_), .A2(new_n599_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n752_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n354_), .B(new_n769_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n758_), .A2(new_n598_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n767_), .B1(new_n778_), .B2(new_n642_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n766_), .B1(new_n779_), .B2(KEYINPUT57), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n767_), .B(new_n781_), .C1(new_n778_), .C2(new_n642_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n324_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n688_), .A2(new_n361_), .A3(new_n360_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT115), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n610_), .A2(new_n786_), .A3(new_n688_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n293_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(new_n293_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n746_), .B1(new_n783_), .B2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n790_), .A2(new_n791_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n752_), .A2(new_n770_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n768_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n773_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n777_), .B1(new_n797_), .B2(KEYINPUT117), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n642_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT57), .B1(new_n800_), .B2(KEYINPUT118), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n289_), .A2(new_n292_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n782_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n612_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n794_), .A2(new_n804_), .A3(KEYINPUT119), .ZN(new_n805_));
  INV_X1    g604(.A(new_n605_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n580_), .A2(new_n806_), .A3(new_n629_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n793_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n599_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n803_), .A2(new_n812_), .A3(new_n612_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n803_), .B2(new_n612_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n794_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n580_), .A2(new_n806_), .A3(KEYINPUT59), .A4(new_n629_), .ZN(new_n816_));
  AOI221_X4 g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .C1(new_n808_), .C2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n808_), .A2(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n816_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n599_), .A2(G113gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n810_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  AND3_X1   g622(.A1(new_n818_), .A2(new_n363_), .A3(new_n819_), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT60), .B2(new_n825_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n824_), .A2(new_n825_), .B1(new_n808_), .B2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n809_), .B2(new_n324_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n324_), .A2(G127gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n821_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n809_), .B2(new_n642_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n650_), .A2(G134gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n821_), .B2(new_n833_), .ZN(G1343gat));
  AND2_X1   g633(.A1(new_n793_), .A2(new_n805_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n806_), .A2(new_n620_), .A3(new_n561_), .A4(new_n579_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n599_), .A3(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n836_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n364_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT122), .B(G148gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1345gat));
  NAND4_X1  g641(.A1(new_n793_), .A2(new_n805_), .A3(new_n324_), .A4(new_n836_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n844_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n839_), .B2(new_n293_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n287_), .A2(G162gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n839_), .B2(new_n852_), .ZN(G1347gat));
  NAND2_X1  g652(.A1(new_n783_), .A2(new_n812_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n814_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n792_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n605_), .A2(new_n568_), .A3(new_n629_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n636_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n693_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT124), .B1(new_n856_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n815_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(G169gat), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n815_), .A2(new_n434_), .A3(new_n861_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n863_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n865_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(G1348gat));
  NOR2_X1   g670(.A1(new_n856_), .A2(new_n860_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G176gat), .B1(new_n872_), .B2(new_n362_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n835_), .A2(new_n561_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n858_), .A2(new_n364_), .A3(new_n428_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1349gat));
  NOR2_X1   g676(.A1(new_n612_), .A2(new_n463_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n872_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT125), .ZN(new_n880_));
  INV_X1    g679(.A(G183gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n857_), .A2(new_n324_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n874_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n879_), .A2(KEYINPUT125), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n872_), .A2(new_n642_), .A3(new_n419_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n872_), .A2(new_n650_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT126), .B1(new_n888_), .B2(G190gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  INV_X1    g689(.A(G190gat), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n890_), .B(new_n891_), .C1(new_n872_), .C2(new_n650_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n887_), .B1(new_n889_), .B2(new_n892_), .ZN(G1351gat));
  AND3_X1   g692(.A1(new_n620_), .A2(new_n562_), .A3(new_n629_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n835_), .A2(new_n599_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n835_), .A2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n364_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n445_), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n835_), .A2(new_n324_), .A3(new_n894_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  OAI21_X1  g703(.A(G218gat), .B1(new_n897_), .B2(new_n293_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n287_), .A2(G218gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n897_), .B2(new_n906_), .ZN(G1355gat));
endmodule


