//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1002_, new_n1003_, new_n1004_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT72), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT70), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(KEYINPUT70), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(KEYINPUT70), .ZN(new_n216_));
  INV_X1    g015(.A(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT15), .A3(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT66), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NOR4_X1   g029(.A1(new_n230_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G85gat), .B(G92gat), .Z(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(KEYINPUT66), .B2(new_n221_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n223_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G85gat), .B(G92gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(KEYINPUT8), .ZN(new_n241_));
  NOR3_X1   g040(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT65), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n222_), .B(new_n241_), .C1(new_n243_), .C2(new_n229_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G85gat), .A2(G92gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT9), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(KEYINPUT9), .B2(new_n239_), .ZN(new_n251_));
  OR2_X1    g050(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n226_), .A3(new_n227_), .A4(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n245_), .B1(new_n251_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT64), .B1(new_n246_), .B2(new_n247_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n236_), .B2(new_n247_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n226_), .A2(new_n227_), .A3(new_n256_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(KEYINPUT67), .A3(new_n255_), .A4(new_n261_), .ZN(new_n262_));
  AND4_X1   g061(.A1(new_n238_), .A2(new_n244_), .A3(new_n258_), .A4(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT71), .B1(new_n220_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G232gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT34), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT35), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n213_), .A2(new_n214_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n260_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n238_), .A2(new_n244_), .A3(new_n271_), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n220_), .A2(new_n263_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n266_), .A2(KEYINPUT35), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n206_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n274_), .B(KEYINPUT73), .C1(new_n273_), .C2(new_n276_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n279_), .A2(new_n280_), .B1(new_n281_), .B2(new_n277_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT25), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n284_), .A2(new_n285_), .B1(KEYINPUT26), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n287_), .B(new_n289_), .C1(new_n285_), .C2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(new_n292_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT82), .B(G176gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n304_), .A2(new_n305_), .B1(G169gat), .B2(G176gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n297_), .B(new_n298_), .C1(G183gat), .C2(G190gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n291_), .A2(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT30), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G71gat), .B(G99gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G43gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G15gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n291_), .A2(new_n303_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n306_), .A2(new_n307_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT30), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n323_), .A2(new_n311_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n318_), .B1(new_n324_), .B2(new_n317_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G134gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G127gat), .ZN(new_n329_));
  INV_X1    g128(.A(G127gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G134gat), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n329_), .A2(new_n331_), .A3(KEYINPUT84), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT84), .B1(new_n329_), .B2(new_n331_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n327_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n331_), .A3(KEYINPUT84), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n326_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n325_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G211gat), .B(G218gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n348_), .A2(new_n349_), .A3(G197gat), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  INV_X1    g150(.A(G204gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT21), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(G197gat), .B1(new_n348_), .B2(new_n349_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT21), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT93), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  OR2_X1    g159(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n351_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n356_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(G218gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G211gat), .ZN(new_n367_));
  INV_X1    g166(.A(G211gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G218gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n351_), .A3(new_n362_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n360_), .B1(G197gat), .B2(G204gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n364_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n355_), .A2(new_n370_), .A3(KEYINPUT21), .A4(new_n357_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT94), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n347_), .A2(new_n360_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n357_), .A4(new_n355_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n359_), .A2(new_n374_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT89), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT88), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n394_));
  NOR4_X1   g193(.A1(new_n394_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n386_), .B(new_n391_), .C1(new_n393_), .C2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n400_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT1), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n399_), .A2(new_n410_), .A3(new_n400_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n411_), .A3(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n387_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n381_), .B1(new_n406_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n380_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n376_), .A2(new_n379_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n354_), .A2(new_n358_), .A3(KEYINPUT93), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n365_), .B1(new_n364_), .B2(new_n373_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n389_), .A2(new_n390_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n392_), .B(KEYINPUT88), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n404_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n415_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n402_), .B1(new_n401_), .B2(KEYINPUT1), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n411_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT29), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n418_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n346_), .B1(new_n420_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT96), .B(new_n346_), .C1(new_n420_), .C2(new_n433_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n419_), .B1(new_n380_), .B2(new_n417_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(new_n432_), .A3(new_n418_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n346_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT95), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n439_), .A3(new_n443_), .A4(new_n440_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n436_), .A2(new_n437_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n446_));
  AOI22_X1  g245(.A1(new_n396_), .A2(new_n405_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT90), .A3(new_n381_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT90), .B1(new_n447_), .B2(new_n381_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n446_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G22gat), .B(G50gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n445_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n458_), .A2(new_n459_), .A3(new_n434_), .A4(new_n441_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT98), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n288_), .A2(G190gat), .ZN(new_n469_));
  INV_X1    g268(.A(G190gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(KEYINPUT26), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n468_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(KEYINPUT26), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n288_), .A2(G190gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT98), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n302_), .B1(new_n476_), .B2(new_n290_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT99), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n299_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n294_), .A2(KEYINPUT99), .A3(new_n297_), .A4(new_n298_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n477_), .A2(new_n481_), .B1(new_n307_), .B2(new_n306_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT20), .B1(new_n380_), .B2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n421_), .B(new_n308_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n467_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n380_), .B2(new_n482_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n424_), .A2(new_n321_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n466_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G8gat), .B(G36gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT18), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n486_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n475_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT98), .B1(new_n473_), .B2(new_n474_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n290_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n302_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n479_), .A2(new_n480_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n320_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT20), .B1(new_n424_), .B2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n380_), .A2(new_n308_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n467_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n487_), .B1(new_n424_), .B2(new_n503_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n466_), .A3(new_n484_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n496_), .B1(new_n509_), .B2(new_n495_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n406_), .A2(new_n416_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n511_), .A2(KEYINPUT101), .A3(KEYINPUT4), .A4(new_n340_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n334_), .A2(new_n339_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT101), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n447_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n447_), .B2(new_n515_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n512_), .B(new_n514_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n340_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n447_), .A2(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n513_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G1gat), .B(G29gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G85gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT0), .B(G57gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n510_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(new_n530_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT33), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n521_), .A2(new_n522_), .A3(new_n514_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n529_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n517_), .A2(new_n519_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n512_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n513_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT102), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n519_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n511_), .A2(KEYINPUT101), .A3(new_n340_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n514_), .B1(new_n548_), .B2(new_n512_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT102), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n536_), .A2(new_n538_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n486_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n494_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT100), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n494_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n504_), .A2(new_n505_), .A3(new_n467_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n466_), .B1(new_n507_), .B2(new_n484_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT100), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n486_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n554_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT103), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n534_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n551_), .A2(KEYINPUT103), .A3(new_n554_), .A4(new_n561_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n463_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n531_), .A2(new_n532_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT27), .B1(new_n558_), .B2(new_n560_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n486_), .A2(new_n490_), .A3(KEYINPUT104), .A4(new_n494_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT104), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n560_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n494_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n570_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n569_), .B1(new_n574_), .B2(KEYINPUT27), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n345_), .B1(new_n566_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n463_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n343_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n533_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n282_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT106), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT11), .ZN(new_n588_));
  XOR2_X1   g387(.A(G71gat), .B(G78gat), .Z(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(KEYINPUT11), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n589_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  INV_X1    g398(.A(G8gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT14), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G1gat), .B(G8gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  AND2_X1   g403(.A1(new_n597_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n597_), .A2(new_n604_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XOR2_X1   g408(.A(G183gat), .B(G211gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n605_), .A2(new_n606_), .B1(new_n607_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n597_), .B(new_n604_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n238_), .A2(new_n244_), .A3(new_n258_), .A4(new_n262_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT68), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n590_), .B(KEYINPUT12), .C1(new_n591_), .C2(new_n592_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n593_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n272_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT12), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n272_), .A2(new_n626_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(new_n625_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n627_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n629_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n625_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT5), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n631_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n631_), .B2(new_n635_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT13), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(KEYINPUT69), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n604_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n215_), .A2(new_n650_), .A3(new_n219_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n218_), .A2(new_n212_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(KEYINPUT76), .A3(new_n604_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT76), .B1(new_n653_), .B2(new_n604_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n651_), .B(new_n652_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT77), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n218_), .A3(new_n212_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n652_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n657_), .A2(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT79), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G169gat), .B(G197gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT78), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n653_), .A2(new_n604_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT76), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n654_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(KEYINPUT77), .A3(new_n652_), .A4(new_n651_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n662_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n668_), .B1(new_n662_), .B2(new_n673_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n649_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n617_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n586_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n567_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n554_), .A2(new_n561_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n532_), .A2(new_n537_), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT33), .B(new_n529_), .C1(new_n520_), .C2(new_n524_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n540_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n549_), .B2(KEYINPUT102), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n543_), .A2(new_n544_), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n684_), .A2(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n563_), .B1(new_n683_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n534_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n565_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n463_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n576_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n343_), .B(KEYINPUT86), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n581_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n677_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(new_n677_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n649_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n277_), .A2(new_n281_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT37), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n277_), .A2(new_n206_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(KEYINPUT37), .B2(new_n282_), .ZN(new_n706_));
  NOR4_X1   g505(.A1(new_n700_), .A2(new_n701_), .A3(new_n617_), .A4(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n599_), .A3(new_n567_), .ZN(new_n708_));
  AOI22_X1  g507(.A1(new_n681_), .A2(G1gat), .B1(new_n682_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n682_), .B2(new_n708_), .ZN(G1324gat));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n600_), .A3(new_n578_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n578_), .B(new_n679_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT39), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(G8gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n712_), .B2(G8gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT40), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(G1325gat));
  NAND3_X1  g517(.A1(new_n707_), .A2(new_n315_), .A3(new_n695_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n680_), .A2(new_n695_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n720_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT41), .B1(new_n720_), .B2(G15gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1326gat));
  INV_X1    g522(.A(G22gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n707_), .A2(new_n724_), .A3(new_n463_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n680_), .A2(new_n463_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G22gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT42), .B(new_n724_), .C1(new_n680_), .C2(new_n463_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1327gat));
  INV_X1    g529(.A(new_n700_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n615_), .B(KEYINPUT75), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n279_), .A2(new_n280_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n702_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n617_), .A2(new_n736_), .A3(new_n282_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n701_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n731_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G29gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n567_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n732_), .A2(new_n678_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT37), .B1(new_n733_), .B2(new_n702_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n703_), .A2(new_n704_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n705_), .B(KEYINPUT107), .C1(KEYINPUT37), .C2(new_n282_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n743_), .B1(new_n696_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n706_), .A2(new_n743_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n742_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT44), .B(new_n742_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G29gat), .B1(new_n757_), .B2(new_n533_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n741_), .A2(new_n758_), .ZN(G1328gat));
  XNOR2_X1  g558(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n575_), .A2(G36gat), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n738_), .B(new_n762_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G36gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n755_), .A2(new_n578_), .A3(new_n756_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(KEYINPUT109), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n755_), .A2(new_n769_), .A3(new_n578_), .A4(new_n756_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n761_), .B(new_n765_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(KEYINPUT109), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(G36gat), .A3(new_n770_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n765_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n760_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n771_), .A2(new_n775_), .ZN(G1329gat));
  INV_X1    g575(.A(new_n757_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(G43gat), .A3(new_n580_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n731_), .A2(new_n695_), .A3(new_n738_), .ZN(new_n779_));
  INV_X1    g578(.A(G43gat), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n779_), .B2(new_n780_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT47), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT47), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n778_), .B(new_n785_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1330gat));
  AOI21_X1  g586(.A(G50gat), .B1(new_n739_), .B2(new_n463_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n463_), .A2(G50gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n777_), .B2(new_n789_), .ZN(G1331gat));
  AOI21_X1  g589(.A(new_n677_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n617_), .A2(new_n706_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n701_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G57gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n567_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n701_), .A2(new_n676_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n617_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n586_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n567_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n800_), .B2(new_n794_), .ZN(G1332gat));
  INV_X1    g600(.A(G64gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n793_), .A2(new_n802_), .A3(new_n578_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n798_), .A2(new_n578_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G64gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT48), .B(new_n802_), .C1(new_n798_), .C2(new_n578_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(G1333gat));
  INV_X1    g607(.A(G71gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n793_), .A2(new_n809_), .A3(new_n695_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n798_), .A2(new_n695_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(G71gat), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G71gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(G1334gat));
  INV_X1    g614(.A(G78gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n793_), .A2(new_n816_), .A3(new_n463_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n463_), .B(new_n797_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(G78gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n818_), .B2(G78gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT113), .ZN(G1335gat));
  AOI21_X1  g622(.A(new_n649_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n791_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G85gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n567_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n750_), .A2(new_n752_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n796_), .A2(new_n732_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n567_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n831_), .B2(new_n826_), .ZN(G1336gat));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n829_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G92gat), .B1(new_n833_), .B2(new_n575_), .ZN(new_n834_));
  INV_X1    g633(.A(G92gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n825_), .A2(new_n835_), .A3(new_n578_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT114), .Z(G1337gat));
  OAI21_X1  g637(.A(G99gat), .B1(new_n833_), .B2(new_n345_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n825_), .A2(new_n580_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g641(.A1(new_n825_), .A2(new_n253_), .A3(new_n463_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n828_), .A2(new_n463_), .A3(new_n829_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(G106gat), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n844_), .B2(G106gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n651_), .B(new_n661_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n666_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n661_), .B1(new_n672_), .B2(new_n659_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n660_), .A2(new_n652_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(KEYINPUT118), .A3(new_n666_), .A4(new_n851_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n662_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n644_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT68), .B1(new_n263_), .B2(new_n620_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n629_), .A2(new_n628_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n632_), .A4(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n865_), .B2(new_n634_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n634_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n624_), .A2(KEYINPUT55), .A3(new_n630_), .A4(new_n625_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n639_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n625_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n631_), .B1(new_n875_), .B2(new_n861_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n640_), .B1(new_n876_), .B2(new_n869_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT56), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n873_), .A2(new_n874_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n641_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n872_), .B(new_n640_), .C1(new_n876_), .C2(new_n869_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(KEYINPUT116), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n860_), .B1(new_n883_), .B2(KEYINPUT117), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n879_), .A2(new_n882_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n282_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n857_), .A2(new_n641_), .A3(new_n858_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT120), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n857_), .A2(new_n890_), .A3(new_n641_), .A4(new_n858_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n873_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n892_), .B(KEYINPUT58), .C1(new_n893_), .C2(new_n881_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n706_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n893_), .B2(new_n881_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n887_), .A2(KEYINPUT57), .B1(new_n894_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n879_), .A2(new_n882_), .A3(new_n885_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n885_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n860_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n903_), .B2(new_n282_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n617_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n792_), .A2(new_n676_), .A3(new_n649_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT54), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n792_), .A2(new_n909_), .A3(new_n676_), .A4(new_n649_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n579_), .A2(new_n567_), .A3(new_n580_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(KEYINPUT59), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n911_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n887_), .B2(KEYINPUT57), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(new_n900_), .C1(new_n903_), .C2(new_n282_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n899_), .A2(new_n917_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n916_), .B1(new_n920_), .B2(new_n617_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n913_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n677_), .B(new_n915_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G113gat), .ZN(new_n925_));
  INV_X1    g724(.A(G113gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n922_), .A2(new_n926_), .A3(new_n677_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1340gat));
  OAI211_X1 g727(.A(new_n701_), .B(new_n915_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G120gat), .ZN(new_n930_));
  INV_X1    g729(.A(G120gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(new_n649_), .B2(KEYINPUT60), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n922_), .B(new_n932_), .C1(KEYINPUT60), .C2(new_n931_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n930_), .A2(new_n933_), .ZN(G1341gat));
  OAI211_X1 g733(.A(new_n732_), .B(new_n915_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G127gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n922_), .A2(new_n330_), .A3(new_n732_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1342gat));
  NAND2_X1  g737(.A1(new_n922_), .A2(new_n282_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n328_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT121), .B(G134gat), .Z(new_n941_));
  NOR2_X1   g740(.A1(new_n895_), .A2(new_n941_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n915_), .B(new_n942_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n940_), .A2(new_n943_), .ZN(G1343gat));
  NAND4_X1  g743(.A1(new_n345_), .A2(new_n567_), .A3(new_n463_), .A4(new_n575_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n921_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n677_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n701_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT122), .B(G148gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1345gat));
  NAND2_X1  g750(.A1(new_n946_), .A2(new_n732_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT61), .B(G155gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1346gat));
  AOI21_X1  g753(.A(G162gat), .B1(new_n946_), .B2(new_n282_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n749_), .A2(G162gat), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n946_), .B2(new_n956_), .ZN(G1347gat));
  NOR3_X1   g756(.A1(new_n345_), .A2(new_n567_), .A3(new_n575_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n732_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n693_), .B(new_n958_), .C1(new_n959_), .C2(new_n916_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G169gat), .B1(new_n960_), .B2(new_n676_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  OAI211_X1 g762(.A(KEYINPUT62), .B(G169gat), .C1(new_n960_), .C2(new_n676_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n463_), .B1(new_n906_), .B2(new_n911_), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n965_), .A2(new_n305_), .A3(new_n677_), .A4(new_n958_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n963_), .A2(new_n964_), .A3(new_n966_), .ZN(G1348gat));
  OAI21_X1  g766(.A(new_n304_), .B1(new_n960_), .B2(new_n649_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(KEYINPUT123), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n970_), .B(new_n304_), .C1(new_n960_), .C2(new_n649_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n921_), .A2(new_n463_), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n958_), .A2(G176gat), .A3(new_n701_), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n969_), .A2(new_n971_), .B1(new_n972_), .B2(new_n973_), .ZN(G1349gat));
  NAND3_X1  g773(.A1(new_n972_), .A2(new_n732_), .A3(new_n958_), .ZN(new_n975_));
  INV_X1    g774(.A(G183gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n958_), .A2(new_n732_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n977_), .A2(new_n290_), .ZN(new_n978_));
  AOI22_X1  g777(.A1(new_n975_), .A2(new_n976_), .B1(new_n965_), .B2(new_n978_), .ZN(G1350gat));
  NAND2_X1  g778(.A1(new_n282_), .A2(new_n476_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n965_), .A2(new_n958_), .A3(new_n981_), .ZN(new_n982_));
  OAI21_X1  g781(.A(G190gat), .B1(new_n960_), .B2(new_n895_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n982_), .A2(new_n983_), .A3(KEYINPUT124), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1351gat));
  NAND3_X1  g787(.A1(new_n345_), .A2(new_n568_), .A3(new_n578_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n920_), .A2(new_n617_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n911_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n677_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n361_), .A2(new_n362_), .ZN(new_n995_));
  INV_X1    g794(.A(new_n995_), .ZN(new_n996_));
  AND4_X1   g795(.A1(new_n994_), .A2(new_n991_), .A3(new_n996_), .A4(new_n701_), .ZN(new_n997_));
  NOR3_X1   g796(.A1(new_n921_), .A2(new_n649_), .A3(new_n989_), .ZN(new_n998_));
  OR2_X1    g797(.A1(new_n998_), .A2(new_n352_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n994_), .B1(new_n998_), .B2(new_n996_), .ZN(new_n1000_));
  AOI21_X1  g799(.A(new_n997_), .B1(new_n999_), .B2(new_n1000_), .ZN(G1353gat));
  AOI21_X1  g800(.A(new_n617_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n991_), .A2(new_n1002_), .ZN(new_n1003_));
  OR2_X1    g802(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1004_));
  XNOR2_X1  g803(.A(new_n1003_), .B(new_n1004_), .ZN(G1354gat));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n1006_));
  AOI21_X1  g805(.A(new_n366_), .B1(new_n991_), .B2(new_n706_), .ZN(new_n1007_));
  NOR4_X1   g806(.A1(new_n921_), .A2(G218gat), .A3(new_n734_), .A4(new_n989_), .ZN(new_n1008_));
  OAI21_X1  g807(.A(new_n1006_), .B1(new_n1007_), .B2(new_n1008_), .ZN(new_n1009_));
  NAND3_X1  g808(.A1(new_n991_), .A2(new_n366_), .A3(new_n282_), .ZN(new_n1010_));
  NOR3_X1   g809(.A1(new_n921_), .A2(new_n895_), .A3(new_n989_), .ZN(new_n1011_));
  OAI211_X1 g810(.A(new_n1010_), .B(KEYINPUT126), .C1(new_n1011_), .C2(new_n366_), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1009_), .A2(new_n1012_), .ZN(G1355gat));
endmodule


