//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT19), .Z(new_n209_));
  OR2_X1    g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(KEYINPUT21), .A3(new_n211_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n215_), .A2(new_n216_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT22), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT93), .Z(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT23), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n235_), .B2(KEYINPUT23), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  INV_X1    g039(.A(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT95), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n232_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(KEYINPUT23), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n234_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT25), .B(G183gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n229_), .A2(KEYINPUT24), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(new_n250_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT92), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n219_), .B1(new_n247_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT20), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n249_), .B2(new_n242_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT22), .B1(new_n223_), .B2(KEYINPUT83), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT83), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n221_), .A3(G169gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n270_), .A3(new_n220_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n229_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n248_), .A2(new_n234_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n266_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n252_), .B1(new_n257_), .B2(new_n250_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n241_), .B2(KEYINPUT26), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G183gat), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT81), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n276_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n273_), .A2(new_n275_), .B1(new_n286_), .B2(new_n239_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n219_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n265_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n209_), .B1(new_n264_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n222_), .A2(new_n224_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT94), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n230_), .B1(new_n294_), .B2(new_n220_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n239_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n245_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n253_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n262_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n261_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n302_), .A3(new_n288_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n209_), .A2(KEYINPUT20), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n254_), .B(new_n278_), .C1(new_n255_), .C2(new_n277_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(new_n239_), .A3(new_n258_), .A4(new_n252_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n275_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n229_), .B(new_n271_), .C1(new_n274_), .C2(new_n266_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n304_), .B1(new_n309_), .B2(new_n219_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n303_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n207_), .B1(new_n290_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n209_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n288_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT20), .B1(new_n309_), .B2(new_n219_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n207_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n310_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT27), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n287_), .A2(new_n288_), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n303_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT103), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n303_), .A2(KEYINPUT103), .A3(new_n322_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n209_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n314_), .A2(new_n315_), .A3(new_n313_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n207_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(KEYINPUT27), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n320_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT87), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n340_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(KEYINPUT1), .B1(new_n337_), .B2(new_n338_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n344_), .A3(new_n343_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n336_), .A2(new_n359_), .A3(new_n340_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n352_), .A2(new_n346_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n333_), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  AOI22_X1  g169(.A1(new_n348_), .A2(new_n357_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  INV_X1    g171(.A(new_n333_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n369_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n219_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n378_));
  AND2_X1   g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n219_), .B2(KEYINPUT89), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OAI221_X1 g180(.A(new_n219_), .B1(KEYINPUT89), .B2(new_n379_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT90), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT91), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n377_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n382_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n377_), .A2(new_n387_), .A3(new_n386_), .A4(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n332_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n309_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT30), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT31), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n406_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n398_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n398_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n358_), .A2(new_n367_), .A3(new_n398_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT96), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n398_), .B1(new_n358_), .B2(new_n367_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n371_), .A2(KEYINPUT96), .A3(new_n398_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n368_), .A2(new_n415_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT96), .A3(new_n418_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n422_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n417_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n431_));
  NOR4_X1   g230(.A1(new_n371_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n398_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n423_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G57gat), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT99), .ZN(new_n436_));
  INV_X1    g235(.A(G1gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n439_));
  INV_X1    g238(.A(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n438_), .A2(new_n441_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n438_), .B(new_n441_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n423_), .B(new_n446_), .C1(new_n428_), .C2(new_n433_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n413_), .A2(new_n416_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n395_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n392_), .A2(new_n445_), .A3(new_n393_), .A4(new_n447_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n332_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n447_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT4), .B1(new_n421_), .B2(new_n422_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT97), .B1(new_n425_), .B2(KEYINPUT4), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n420_), .A2(new_n430_), .A3(new_n424_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n417_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT33), .A3(new_n423_), .A4(new_n446_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n312_), .A2(new_n319_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n429_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n444_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT100), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n429_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n466_), .A2(new_n467_), .B1(new_n457_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(KEYINPUT100), .A3(new_n444_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n464_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n316_), .A2(new_n318_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n205_), .A2(KEYINPUT32), .A3(new_n206_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT101), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n463_), .A2(new_n471_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n394_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n454_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n413_), .A2(new_n416_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n451_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n484_), .A2(new_n485_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G1gat), .A2(G8gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT14), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n437_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .A4(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n489_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n484_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n486_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n489_), .A2(new_n499_), .A3(KEYINPUT77), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT78), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT78), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n507_), .A2(new_n513_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n508_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n503_), .A2(KEYINPUT15), .A3(new_n486_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n499_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n518_), .A2(KEYINPUT79), .A3(new_n499_), .A4(new_n519_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n516_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n515_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT80), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n515_), .B2(new_n525_), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n530_), .B(new_n524_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n483_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  OAI22_X1  g340(.A1(new_n541_), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n541_), .B2(KEYINPUT9), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT66), .B(G92gat), .ZN(new_n544_));
  INV_X1    g343(.A(G85gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n540_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G106gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT64), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n548_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT6), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n547_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  OR4_X1    g356(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  INV_X1    g358(.A(G99gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n548_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT7), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n564_));
  XOR2_X1   g363(.A(G85gat), .B(G92gat), .Z(new_n565_));
  AND3_X1   g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n557_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n570_));
  XOR2_X1   g369(.A(G71gat), .B(G78gat), .Z(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n557_), .B(new_n575_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT12), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n568_), .A2(new_n580_), .A3(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n583_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n590_), .B1(new_n594_), .B2(new_n585_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n592_), .A2(KEYINPUT69), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT69), .B1(new_n592_), .B2(new_n595_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT13), .ZN(new_n599_));
  AND2_X1   g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n575_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT75), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n601_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n499_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT76), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n603_), .A2(new_n606_), .A3(new_n607_), .A4(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n603_), .A2(new_n606_), .A3(new_n612_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT76), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT72), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT73), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n568_), .A2(new_n519_), .A3(new_n518_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n557_), .B(new_n504_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT35), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n628_), .A2(new_n637_), .A3(new_n633_), .A4(new_n634_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n627_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n623_), .B(KEYINPUT36), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT74), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT37), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT74), .B(KEYINPUT37), .C1(new_n639_), .C2(new_n642_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n620_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n539_), .A2(new_n599_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n437_), .A3(new_n448_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT104), .Z(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n652_));
  INV_X1    g451(.A(new_n538_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n599_), .A2(new_n653_), .A3(new_n620_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT105), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n639_), .A2(new_n642_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n483_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(KEYINPUT105), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n449_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n651_), .A2(new_n652_), .A3(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n332_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n494_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n659_), .B2(new_n332_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n663_), .B(new_n664_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n665_), .B(KEYINPUT39), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n664_), .B1(new_n670_), .B2(new_n663_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n659_), .B2(new_n482_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n482_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n648_), .A2(new_n403_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n659_), .B2(new_n394_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n648_), .A2(new_n685_), .A3(new_n480_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n620_), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n539_), .A2(new_n599_), .A3(new_n688_), .A4(new_n656_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n440_), .A3(new_n448_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n599_), .A2(new_n653_), .A3(new_n688_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n645_), .A2(new_n646_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n483_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n477_), .A2(new_n478_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n464_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n417_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n467_), .B1(new_n697_), .B2(new_n446_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n457_), .A2(new_n468_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n470_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n696_), .A2(new_n700_), .A3(new_n456_), .A4(new_n462_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n480_), .B1(new_n695_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n328_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n303_), .A2(KEYINPUT103), .A3(new_n322_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT103), .B1(new_n303_), .B2(new_n322_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n321_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n706_), .B2(new_n209_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n330_), .B1(new_n707_), .B2(new_n207_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n452_), .A3(new_n320_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n482_), .B1(new_n702_), .B2(new_n709_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n395_), .A2(new_n450_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n645_), .A2(new_n646_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n692_), .B1(new_n694_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n448_), .B1(new_n716_), .B2(KEYINPUT44), .ZN(new_n717_));
  INV_X1    g516(.A(new_n692_), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT43), .B(new_n693_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n713_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n718_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT108), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n723_), .A3(KEYINPUT44), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n717_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n440_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n722_), .A2(new_n724_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n449_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n726_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n691_), .B1(new_n727_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n721_), .A2(KEYINPUT108), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n723_), .B1(new_n716_), .B2(KEYINPUT44), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n726_), .B(new_n731_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G29gat), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(KEYINPUT110), .A3(new_n732_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n690_), .B1(new_n734_), .B2(new_n739_), .ZN(G1328gat));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n332_), .A2(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n332_), .A2(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n689_), .A2(new_n741_), .A3(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT45), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n332_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n747_), .B(new_n748_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G36gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n728_), .B2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT46), .B(new_n746_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1329gat));
  NAND2_X1  g555(.A1(new_n729_), .A2(new_n730_), .ZN(new_n757_));
  AND4_X1   g556(.A1(G43gat), .A2(new_n728_), .A3(new_n676_), .A4(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G43gat), .B1(new_n689_), .B2(new_n676_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n758_), .A2(KEYINPUT47), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT47), .B1(new_n758_), .B2(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n689_), .B2(new_n480_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n728_), .A2(new_n757_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n480_), .A2(G50gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1331gat));
  NOR3_X1   g565(.A1(new_n599_), .A2(new_n653_), .A3(new_n688_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n657_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n449_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n599_), .A2(new_n653_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n712_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n688_), .A3(new_n714_), .ZN(new_n773_));
  INV_X1    g572(.A(G57gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n448_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(G1332gat));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(new_n744_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n744_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G64gat), .B1(new_n769_), .B2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT48), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT48), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT113), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n768_), .B2(new_n676_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT49), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n773_), .A2(new_n785_), .A3(new_n676_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1334gat));
  INV_X1    g588(.A(G78gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n768_), .B2(new_n480_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT50), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n790_), .A3(new_n480_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1335gat));
  INV_X1    g593(.A(new_n656_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n772_), .A2(new_n620_), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n545_), .A3(new_n448_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n771_), .A2(new_n688_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n694_), .B2(new_n715_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(new_n448_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n800_), .B2(new_n545_), .ZN(G1336gat));
  AOI21_X1  g600(.A(G92gat), .B1(new_n796_), .B2(new_n662_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n779_), .A2(new_n544_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n799_), .B2(new_n803_), .ZN(G1337gat));
  AOI21_X1  g603(.A(new_n560_), .B1(new_n799_), .B2(new_n676_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n552_), .A2(new_n553_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n482_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n796_), .B2(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g608(.A1(new_n796_), .A2(new_n548_), .A3(new_n480_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n799_), .A2(new_n480_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G106gat), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT52), .B(new_n548_), .C1(new_n799_), .C2(new_n480_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g615(.A1(new_n395_), .A2(new_n449_), .A3(new_n482_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n533_), .A2(new_n537_), .A3(new_n592_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n579_), .A2(new_n593_), .A3(new_n581_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n584_), .A2(KEYINPUT55), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n591_), .B1(new_n594_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT115), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n522_), .A2(new_n523_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n509_), .A3(new_n505_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n530_), .A3(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n532_), .A2(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n827_), .A2(new_n832_), .B1(new_n598_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n819_), .B1(new_n838_), .B2(new_n656_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n597_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n592_), .A2(KEYINPUT69), .A3(new_n595_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n837_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n821_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n579_), .A2(new_n593_), .A3(new_n581_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(new_n594_), .A3(new_n824_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n582_), .A2(new_n824_), .A3(new_n583_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n590_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n848_), .A2(new_n533_), .A3(new_n537_), .A4(new_n592_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n829_), .B2(KEYINPUT115), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n842_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n795_), .A3(KEYINPUT57), .ZN(new_n852_));
  NOR2_X1   g651(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n823_), .B(new_n825_), .C1(KEYINPUT116), .C2(KEYINPUT56), .ZN(new_n855_));
  NAND2_X1  g654(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n837_), .A2(new_n592_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(KEYINPUT58), .A3(new_n858_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n714_), .A3(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n839_), .A2(new_n852_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT117), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n839_), .A2(new_n863_), .A3(new_n866_), .A4(new_n852_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n688_), .A3(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n598_), .A2(KEYINPUT13), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n598_), .A2(KEYINPUT13), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n647_), .B(new_n538_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n818_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G113gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n653_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n864_), .A2(new_n688_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n873_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n818_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT118), .B1(new_n875_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n620_), .B1(new_n864_), .B2(KEYINPUT117), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n873_), .B1(new_n884_), .B2(new_n867_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n883_), .B(KEYINPUT59), .C1(new_n885_), .C2(new_n818_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n538_), .B(new_n880_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n877_), .B1(new_n887_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n599_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n875_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n599_), .B(new_n880_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g692(.A(G127gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n875_), .A2(new_n894_), .A3(new_n620_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n688_), .B(new_n880_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1342gat));
  INV_X1    g696(.A(G134gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n875_), .A2(new_n898_), .A3(new_n656_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n693_), .B(new_n880_), .C1(new_n882_), .C2(new_n886_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1343gat));
  NOR4_X1   g700(.A1(new_n744_), .A2(new_n394_), .A3(new_n449_), .A4(new_n676_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n885_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n653_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n868_), .A2(new_n874_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n653_), .A3(new_n902_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT120), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT119), .B(G141gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1344gat));
  INV_X1    g711(.A(new_n599_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n904_), .A2(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n904_), .A2(KEYINPUT121), .A3(new_n620_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n907_), .A2(new_n620_), .A3(new_n902_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  NAND2_X1  g721(.A1(new_n907_), .A2(new_n902_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n693_), .ZN(new_n924_));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n656_), .A2(new_n925_), .ZN(new_n926_));
  OAI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929_));
  OAI221_X1 g728(.A(new_n929_), .B1(new_n923_), .B2(new_n926_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n779_), .A2(new_n450_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n394_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n879_), .A2(new_n933_), .ZN(new_n934_));
  AOI211_X1 g733(.A(KEYINPUT62), .B(new_n223_), .C1(new_n934_), .C2(new_n653_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n653_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(G169gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n934_), .A2(new_n653_), .A3(new_n294_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1348gat));
  AOI21_X1  g739(.A(G176gat), .B1(new_n934_), .B2(new_n913_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n885_), .B2(new_n480_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n907_), .A2(KEYINPUT123), .A3(new_n394_), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n943_), .A2(new_n944_), .A3(new_n932_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n599_), .A2(new_n220_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n941_), .B1(new_n945_), .B2(new_n946_), .ZN(G1349gat));
  INV_X1    g746(.A(new_n934_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n948_), .A2(new_n254_), .A3(new_n688_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n945_), .A2(new_n620_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n240_), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n948_), .B2(new_n693_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n934_), .A2(new_n255_), .A3(new_n656_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1351gat));
  NAND2_X1  g753(.A1(new_n482_), .A2(new_n453_), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n955_), .B(KEYINPUT124), .Z(new_n956_));
  NOR3_X1   g755(.A1(new_n885_), .A2(new_n779_), .A3(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n653_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g758(.A(G204gat), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n957_), .B(new_n913_), .C1(KEYINPUT125), .C2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(KEYINPUT125), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(KEYINPUT126), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n961_), .B(new_n963_), .ZN(G1353gat));
  NAND2_X1  g763(.A1(new_n957_), .A2(new_n620_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(KEYINPUT63), .B(G211gat), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n965_), .B2(new_n968_), .ZN(G1354gat));
  INV_X1    g768(.A(G218gat), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n957_), .A2(new_n970_), .A3(new_n656_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n957_), .A2(new_n714_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n970_), .ZN(G1355gat));
endmodule


