//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT65), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n207_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G85gat), .B(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n204_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT65), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n214_), .B2(new_n215_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(KEYINPUT66), .B(new_n219_), .C1(new_n224_), .C2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n218_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n210_), .A2(new_n212_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n207_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT9), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n226_), .B2(KEYINPUT9), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT64), .ZN(new_n236_));
  OAI221_X1 g035(.A(new_n234_), .B1(new_n222_), .B2(new_n223_), .C1(new_n236_), .C2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G29gat), .B(G36gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT71), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G43gat), .B(G50gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n239_), .A2(KEYINPUT71), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(KEYINPUT71), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n241_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT35), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT34), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n249_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n238_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n230_), .A2(KEYINPUT67), .A3(new_n237_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(KEYINPUT15), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n243_), .A2(new_n246_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .A4(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n253_), .A2(new_n255_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n255_), .B1(new_n253_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n203_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G190gat), .B(G218gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n269_), .B(new_n203_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n264_), .A2(new_n265_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n202_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n278_));
  AOI211_X1 g077(.A(KEYINPUT37), .B(new_n276_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G127gat), .B(G155gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT16), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G183gat), .B(G211gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT74), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n294_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n284_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n284_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(KEYINPUT17), .B2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(KEYINPUT17), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n280_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT76), .Z(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(G85gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G57gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(G155gat), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT1), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  AND4_X1   g120(.A1(KEYINPUT85), .A2(new_n318_), .A3(new_n319_), .A4(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(new_n321_), .C2(KEYINPUT85), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT87), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT3), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n325_), .B(KEYINPUT2), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n323_), .B2(new_n329_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n332_), .B(new_n333_), .C1(new_n331_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  XOR2_X1   g136(.A(G155gat), .B(G162gat), .Z(new_n338_));
  AND3_X1   g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n328_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT89), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT89), .B(new_n328_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G127gat), .B(G134gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n341_), .A2(new_n347_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n354_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n315_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n353_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(G225gat), .A3(G233gat), .A4(new_n350_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n315_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n363_), .A3(KEYINPUT94), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n361_), .A2(new_n365_), .A3(new_n362_), .A4(new_n357_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(G197gat), .ZN(new_n374_));
  INV_X1    g173(.A(G197gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(G204gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT21), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n374_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n379_), .B2(new_n374_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n377_), .B(new_n378_), .C1(new_n381_), .C2(KEYINPUT21), .ZN(new_n382_));
  INV_X1    g181(.A(new_n378_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(KEYINPUT21), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT23), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(G183gat), .A3(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G169gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G169gat), .ZN(new_n395_));
  INV_X1    g194(.A(G176gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT24), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398_));
  MUX2_X1   g197(.A(new_n397_), .B(KEYINPUT24), .S(new_n398_), .Z(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT25), .B(G183gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT82), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(KEYINPUT82), .B2(new_n389_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n394_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n372_), .B1(new_n385_), .B2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409_));
  NAND2_X1  g208(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n408_), .B(KEYINPUT25), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(new_n400_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(KEYINPUT81), .A3(new_n413_), .A4(new_n400_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n390_), .A3(new_n417_), .A4(new_n399_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n408_), .A2(new_n410_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(G190gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n393_), .B1(new_n405_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n407_), .B1(new_n422_), .B2(new_n385_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n426_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n385_), .A2(new_n406_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(new_n372_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(new_n385_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n371_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n423_), .A2(new_n426_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n371_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n438_), .A2(KEYINPUT93), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT93), .B1(new_n438_), .B2(new_n439_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n435_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n364_), .A2(new_n366_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n359_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT33), .B(new_n315_), .C1(new_n355_), .C2(new_n358_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n370_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n436_), .A2(new_n437_), .A3(new_n370_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n354_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n362_), .C1(new_n356_), .C2(new_n354_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n445_), .A2(new_n446_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n443_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G71gat), .B(G99gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G43gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n422_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n418_), .A2(new_n421_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(G15gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT30), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n465_), .A3(new_n460_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n455_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n347_), .B(KEYINPUT31), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n469_), .B2(new_n455_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n455_), .B(new_n473_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G22gat), .B(G50gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n343_), .A2(KEYINPUT29), .A3(new_n344_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT90), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n336_), .A2(new_n338_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT88), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n327_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n385_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n484_), .A2(new_n487_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT29), .B1(new_n343_), .B2(new_n344_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI211_X1 g297(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n343_), .C2(new_n344_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n495_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n483_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n484_), .A2(new_n487_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n494_), .A2(new_n488_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n500_), .A3(new_n482_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n479_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n448_), .A2(new_n449_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(KEYINPUT27), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n447_), .B1(new_n427_), .B2(new_n433_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT95), .B(new_n447_), .C1(new_n427_), .C2(new_n433_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n449_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n519_), .B2(KEYINPUT27), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n509_), .A2(new_n500_), .A3(new_n482_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n482_), .B1(new_n509_), .B2(new_n500_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n479_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n477_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n520_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n364_), .A2(new_n366_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n454_), .A2(new_n512_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n289_), .A2(KEYINPUT12), .A3(new_n290_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n257_), .A2(new_n258_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT68), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n230_), .A2(new_n237_), .A3(new_n291_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n291_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n257_), .A2(new_n538_), .A3(new_n258_), .A4(new_n530_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n536_), .A3(new_n537_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n533_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n534_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G176gat), .B(G204gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT70), .ZN(new_n546_));
  XOR2_X1   g345(.A(G120gat), .B(G148gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n550_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n543_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(KEYINPUT13), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n301_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n259_), .A2(new_n262_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n260_), .A2(new_n301_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n247_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n563_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G113gat), .B(G141gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT77), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n564_), .A2(new_n568_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT78), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n559_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n528_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n311_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n527_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n296_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT38), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n276_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n528_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n577_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n308_), .A2(new_n558_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n527_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(G1324gat));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n297_), .A3(new_n520_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n520_), .A3(new_n589_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(G8gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n594_), .B2(G8gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g399(.A(G15gat), .B1(new_n590_), .B2(new_n479_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n581_), .A2(new_n463_), .A3(new_n524_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1326gat));
  NAND2_X1  g403(.A1(new_n503_), .A2(new_n510_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G22gat), .B1(new_n590_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT42), .ZN(new_n608_));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n581_), .A2(new_n609_), .A3(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(G1327gat));
  NOR2_X1   g410(.A1(KEYINPUT98), .A2(KEYINPUT44), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n309_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n558_), .A2(new_n588_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n617_), .B(KEYINPUT43), .C1(new_n528_), .C2(new_n280_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n278_), .A2(new_n279_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n523_), .A2(new_n525_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n520_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n621_), .A2(new_n527_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n511_), .B1(new_n443_), .B2(new_n453_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT43), .B1(new_n625_), .B2(new_n617_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n616_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT98), .B1(KEYINPUT97), .B2(KEYINPUT44), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n617_), .B1(new_n528_), .B2(new_n280_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n618_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n616_), .A3(new_n628_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n527_), .B1(new_n630_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n309_), .A2(new_n585_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n580_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n582_), .A2(new_n637_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT99), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n636_), .A2(new_n637_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT100), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(KEYINPUT100), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n630_), .A2(new_n635_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n520_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n639_), .A2(G36gat), .A3(new_n622_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n644_), .B(new_n645_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n628_), .B1(new_n634_), .B2(new_n616_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n615_), .B(new_n629_), .C1(new_n633_), .C2(new_n618_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n520_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G36gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n650_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(KEYINPUT100), .A3(new_n656_), .A4(new_n643_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n651_), .A2(new_n657_), .ZN(G1329gat));
  INV_X1    g457(.A(G43gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n647_), .B2(new_n524_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n639_), .A2(G43gat), .A3(new_n479_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1330gat));
  INV_X1    g464(.A(new_n639_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G50gat), .B1(new_n666_), .B2(new_n605_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n605_), .A2(G50gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n647_), .B2(new_n668_), .ZN(G1331gat));
  NOR3_X1   g468(.A1(new_n559_), .A2(new_n308_), .A3(new_n578_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n587_), .A2(new_n582_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G57gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n558_), .A2(new_n588_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n528_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n311_), .A2(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n527_), .A2(G57gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(G1332gat));
  NAND3_X1  g476(.A1(new_n587_), .A2(new_n520_), .A3(new_n670_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT48), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(G64gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n678_), .B2(G64gat), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n622_), .A2(G64gat), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n681_), .A2(new_n682_), .B1(new_n675_), .B2(new_n683_), .ZN(G1333gat));
  NAND3_X1  g483(.A1(new_n587_), .A2(new_n524_), .A3(new_n670_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT101), .B(KEYINPUT49), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(G71gat), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n685_), .B2(G71gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n479_), .A2(G71gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT102), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n688_), .A2(new_n689_), .B1(new_n675_), .B2(new_n691_), .ZN(G1334gat));
  NAND3_X1  g491(.A1(new_n587_), .A2(new_n605_), .A3(new_n670_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT50), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(G78gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n693_), .B2(G78gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n606_), .A2(G78gat), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT103), .Z(new_n699_));
  OAI22_X1  g498(.A1(new_n696_), .A2(new_n697_), .B1(new_n675_), .B2(new_n699_), .ZN(G1335gat));
  NAND2_X1  g499(.A1(new_n674_), .A2(new_n638_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n582_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n634_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n309_), .A2(new_n673_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT104), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT104), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n704_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n582_), .A2(G85gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT105), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n703_), .B1(new_n710_), .B2(new_n712_), .ZN(G1336gat));
  NAND3_X1  g512(.A1(new_n702_), .A2(new_n232_), .A3(new_n520_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n704_), .A2(new_n709_), .A3(new_n622_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n232_), .ZN(G1337gat));
  OR3_X1    g515(.A1(new_n701_), .A2(new_n236_), .A3(new_n479_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n634_), .A2(new_n708_), .A3(new_n524_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT106), .A3(G99gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n718_), .B2(G99gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n634_), .A2(new_n708_), .A3(new_n605_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT52), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT108), .B1(new_n723_), .B2(G106gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n634_), .A2(new_n708_), .A3(new_n605_), .ZN(new_n731_));
  INV_X1    g530(.A(G106gat), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n730_), .B(new_n725_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n702_), .A2(new_n732_), .A3(new_n605_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT53), .B1(new_n729_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n726_), .A3(new_n724_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n733_), .A4(new_n734_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1339gat));
  XNOR2_X1  g540(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n558_), .A2(new_n578_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n310_), .B2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n280_), .A2(new_n309_), .A3(new_n744_), .A4(new_n742_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(KEYINPUT114), .A2(KEYINPUT58), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n561_), .A2(new_n563_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT110), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n561_), .A2(new_n754_), .A3(new_n563_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n753_), .A2(new_n567_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n566_), .A2(new_n562_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n573_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n751_), .B(new_n576_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n562_), .B1(new_n752_), .B2(KEYINPUT110), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n760_), .B2(new_n755_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n576_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT111), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n759_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n553_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n535_), .B1(new_n531_), .B2(KEYINPUT68), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n537_), .B1(new_n766_), .B2(new_n539_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n540_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n766_), .A2(KEYINPUT55), .A3(new_n537_), .A4(new_n539_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n550_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n552_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n765_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n280_), .B1(new_n750_), .B2(new_n775_), .ZN(new_n776_));
  AND4_X1   g575(.A1(new_n537_), .A2(new_n532_), .A3(new_n539_), .A4(new_n536_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n532_), .A2(new_n539_), .A3(new_n536_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n541_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(KEYINPUT55), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n770_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n550_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n773_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n550_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n750_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n765_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n553_), .A2(new_n577_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n764_), .A2(new_n554_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n586_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n776_), .A2(new_n787_), .B1(new_n791_), .B2(KEYINPUT57), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  INV_X1    g594(.A(new_n793_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n790_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n795_), .B(new_n796_), .C1(new_n798_), .C2(new_n586_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n794_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n749_), .B1(new_n800_), .B2(new_n308_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n527_), .A2(new_n520_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n525_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806_), .B2(new_n577_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n791_), .A2(new_n793_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n309_), .B1(new_n792_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n749_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n804_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n799_), .A2(new_n794_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n775_), .A2(new_n750_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n787_), .A2(new_n816_), .A3(new_n620_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n789_), .A2(new_n790_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n585_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n817_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n308_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n748_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n804_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(KEYINPUT59), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n578_), .A2(G113gat), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT115), .Z(new_n827_));
  AOI21_X1  g626(.A(new_n807_), .B1(new_n825_), .B2(new_n827_), .ZN(G1340gat));
  OAI22_X1  g627(.A1(new_n806_), .A2(new_n812_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G120gat), .B1(new_n829_), .B2(new_n559_), .ZN(new_n830_));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n559_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(KEYINPUT60), .B2(new_n831_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n824_), .B2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n806_), .B2(new_n309_), .ZN(new_n835_));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n309_), .B2(KEYINPUT116), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(KEYINPUT116), .B2(new_n836_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n835_), .B1(new_n825_), .B2(new_n838_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n824_), .B2(new_n585_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT117), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n840_), .C1(new_n824_), .C2(new_n585_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n280_), .A2(new_n840_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT118), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n842_), .A2(new_n844_), .B1(new_n825_), .B2(new_n846_), .ZN(G1343gat));
  AOI21_X1  g646(.A(new_n523_), .B1(new_n822_), .B2(new_n748_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n577_), .A3(new_n802_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n558_), .A3(new_n802_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT119), .B(G148gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1345gat));
  INV_X1    g652(.A(new_n523_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n823_), .A2(new_n854_), .A3(new_n309_), .A4(new_n802_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT120), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n848_), .A2(new_n857_), .A3(new_n309_), .A4(new_n802_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n856_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1346gat));
  NAND4_X1  g661(.A1(new_n848_), .A2(new_n317_), .A3(new_n586_), .A4(new_n802_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n801_), .A2(new_n523_), .A3(new_n280_), .A4(new_n803_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n317_), .ZN(G1347gat));
  NAND2_X1  g664(.A1(new_n527_), .A2(new_n520_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n866_), .A2(new_n525_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n811_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT22), .B(G169gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n577_), .A3(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n866_), .A2(new_n479_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n577_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n872_), .A2(KEYINPUT121), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(KEYINPUT121), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n875_), .B(new_n606_), .C1(new_n810_), .C2(new_n749_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(KEYINPUT122), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n877_));
  OR2_X1    g676(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n606_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n308_), .B1(new_n821_), .B2(new_n808_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n748_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n878_), .B(new_n879_), .C1(new_n882_), .C2(new_n395_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n870_), .A2(new_n877_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n870_), .A2(new_n883_), .A3(new_n886_), .A4(new_n877_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n868_), .B2(new_n558_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n801_), .A2(new_n605_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n559_), .A2(new_n866_), .A3(new_n396_), .A4(new_n479_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  INV_X1    g691(.A(new_n868_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(new_n401_), .A3(new_n308_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n419_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n309_), .A3(new_n871_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n893_), .B2(new_n280_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n868_), .A2(new_n586_), .A3(new_n400_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1351gat));
  INV_X1    g699(.A(new_n866_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n848_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n588_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n375_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n559_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n373_), .A2(KEYINPUT124), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n373_), .A2(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n907_), .ZN(G1353gat));
  NOR2_X1   g708(.A1(new_n902_), .A2(new_n308_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(new_n911_), .ZN(G1354gat));
  XNOR2_X1  g713(.A(KEYINPUT125), .B(G218gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n620_), .A2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT126), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n848_), .A2(new_n901_), .A3(new_n917_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n801_), .A2(new_n585_), .A3(new_n523_), .A4(new_n866_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n915_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n922_), .B(new_n918_), .C1(new_n919_), .C2(new_n915_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1355gat));
endmodule


