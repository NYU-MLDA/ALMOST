//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n212_), .B2(KEYINPUT9), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(new_n212_), .B2(KEYINPUT9), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(KEYINPUT65), .A3(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n209_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n203_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n212_), .A2(new_n214_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n224_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G57gat), .B(G64gat), .Z(new_n235_));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G78gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n220_), .A2(new_n222_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n228_), .A2(new_n225_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n231_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n224_), .A3(new_n244_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n202_), .B1(new_n246_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT66), .ZN(new_n255_));
  INV_X1    g054(.A(new_n224_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(KEYINPUT67), .A3(new_n251_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n242_), .A2(new_n261_), .A3(new_n243_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT12), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n260_), .B2(new_n265_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n232_), .A2(new_n233_), .A3(new_n257_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n250_), .B2(new_n251_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n224_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n244_), .A2(KEYINPUT68), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n262_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT12), .B1(new_n234_), .B2(new_n245_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n253_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n266_), .A2(new_n274_), .A3(new_n277_), .A4(new_n202_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n255_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  AND4_X1   g082(.A1(new_n202_), .A2(new_n266_), .A3(new_n274_), .A4(new_n277_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n254_), .B(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n282_), .B(KEYINPUT70), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n283_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT13), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT13), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(new_n283_), .C1(new_n287_), .C2(new_n289_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G29gat), .B(G36gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT71), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306_));
  INV_X1    g105(.A(G22gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(KEYINPUT74), .A2(G15gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT74), .A2(G15gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312_));
  INV_X1    g111(.A(G15gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G22gat), .A3(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT14), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(G1gat), .B2(G8gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n306_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT75), .B(new_n318_), .C1(new_n311_), .C2(new_n315_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G1gat), .B(G8gat), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n309_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n325_));
  AOI21_X1  g124(.A(G22gat), .B1(new_n314_), .B2(new_n308_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n319_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT75), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n316_), .A2(new_n306_), .A3(new_n319_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n305_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n322_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n303_), .A2(new_n304_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(KEYINPUT76), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G229gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n323_), .A2(new_n330_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n334_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n303_), .A2(KEYINPUT15), .A3(new_n304_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT15), .B1(new_n303_), .B2(new_n304_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n333_), .B(new_n332_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n337_), .A3(new_n331_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G141gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G169gat), .B(G197gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT80), .ZN(new_n354_));
  INV_X1    g153(.A(new_n352_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(new_n346_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n347_), .A2(new_n359_), .A3(new_n352_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n357_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n363_));
  AOI211_X1 g162(.A(KEYINPUT80), .B(new_n355_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(G231gat), .A2(G233gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n339_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n262_), .A3(new_n272_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G127gat), .B(G155gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT16), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G183gat), .B(G211gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n369_), .A2(new_n244_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(new_n245_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n375_), .B(KEYINPUT17), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n294_), .A2(new_n366_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT100), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT89), .B(G106gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT3), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(KEYINPUT3), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n393_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n392_), .A2(KEYINPUT1), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n392_), .A2(KEYINPUT1), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n391_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n395_), .A2(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT28), .B1(new_n409_), .B2(KEYINPUT29), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n393_), .A2(new_n402_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G211gat), .B(G218gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT88), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G197gat), .B(G204gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n418_), .A2(new_n419_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n417_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n415_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G22gat), .B(G50gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n424_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(G78gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n431_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n426_), .A2(new_n429_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n427_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n440_), .B2(new_n430_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n388_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n435_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n430_), .A3(new_n437_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n387_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446_));
  INV_X1    g245(.A(G43gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT30), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT22), .ZN(new_n450_));
  OR2_X1    g249(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G176gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT83), .B1(new_n450_), .B2(G169gat), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n455_), .B(new_n456_), .C1(new_n453_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT23), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(G183gat), .B2(G190gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT25), .B(G183gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT26), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT81), .B1(new_n465_), .B2(G190gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT26), .B(G190gat), .Z(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G169gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n456_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT24), .A3(new_n459_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n461_), .B(new_n473_), .C1(KEYINPUT24), .C2(new_n472_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n463_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n463_), .A2(new_n475_), .A3(KEYINPUT84), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G227gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(new_n313_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n449_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n449_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n483_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490_));
  XOR2_X1   g289(.A(G127gat), .B(G134gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G113gat), .B(G120gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT31), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n494_), .B2(KEYINPUT85), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n486_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n486_), .A2(new_n489_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n494_), .A2(new_n490_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n495_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n496_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n442_), .A2(new_n445_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G29gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G57gat), .B(G85gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  OR4_X1    g307(.A1(KEYINPUT94), .A2(new_n411_), .A3(KEYINPUT4), .A4(new_n493_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n510_));
  INV_X1    g309(.A(new_n493_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n409_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n411_), .A2(new_n493_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT4), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n411_), .B(new_n511_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n508_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n507_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n509_), .A2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n508_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n507_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n519_), .A2(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n518_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n521_), .B2(new_n508_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT33), .A4(new_n507_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n424_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n478_), .A2(new_n530_), .A3(new_n479_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n469_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(new_n464_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n474_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n462_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G169gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n456_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n459_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n536_), .A2(KEYINPUT92), .A3(new_n541_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n534_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT20), .B(new_n531_), .C1(new_n546_), .C2(new_n530_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G226gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT19), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G8gat), .B(G36gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G64gat), .B(G92gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n549_), .B1(new_n546_), .B2(new_n530_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n478_), .A2(new_n479_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n424_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n550_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n549_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n531_), .A2(KEYINPUT20), .ZN(new_n564_));
  INV_X1    g363(.A(new_n534_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n545_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT92), .B1(new_n536_), .B2(new_n541_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n424_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n563_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n530_), .B(new_n565_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n560_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n555_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT96), .B1(new_n519_), .B2(new_n520_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n529_), .A2(new_n562_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n526_), .B(new_n507_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n547_), .A2(new_n549_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n555_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n547_), .A2(new_n549_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n530_), .A2(new_n565_), .A3(new_n542_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n563_), .B1(new_n560_), .B2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT32), .B(new_n556_), .C1(new_n580_), .C2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n502_), .B1(new_n575_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT27), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n570_), .A2(new_n572_), .A3(new_n555_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n556_), .B1(new_n550_), .B2(new_n561_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n573_), .A2(new_n562_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT98), .A3(new_n586_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n555_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT27), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT97), .B1(new_n577_), .B2(new_n556_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(KEYINPUT97), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n591_), .A2(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n443_), .A2(new_n444_), .A3(new_n387_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n387_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n501_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n500_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n442_), .A2(new_n445_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n576_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n585_), .B1(new_n599_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n343_), .A2(new_n344_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n260_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n234_), .A2(new_n334_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT35), .B(new_n609_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n269_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(KEYINPUT72), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n613_), .A2(new_n618_), .A3(KEYINPUT72), .A4(new_n623_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n607_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n386_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT101), .Z(new_n634_));
  INV_X1    g433(.A(new_n576_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n524_), .A2(new_n528_), .A3(new_n574_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n584_), .B1(new_n592_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n600_), .A2(new_n601_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n501_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n600_), .A2(new_n601_), .A3(new_n501_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n604_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n635_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n562_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n598_), .A2(KEYINPUT27), .A3(new_n645_), .A4(new_n594_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n592_), .B2(new_n586_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n590_), .B(KEYINPUT27), .C1(new_n573_), .C2(new_n562_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n640_), .B1(new_n643_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n294_), .A2(new_n366_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n627_), .A2(new_n630_), .A3(new_n653_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n383_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n652_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G1gat), .A3(new_n635_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n636_), .A2(new_n662_), .ZN(G1324gat));
  NAND3_X1  g462(.A1(new_n386_), .A2(new_n632_), .A3(new_n649_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT102), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT102), .ZN(new_n666_));
  INV_X1    g465(.A(G8gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(KEYINPUT39), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n666_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT103), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT103), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n665_), .A2(new_n666_), .A3(new_n669_), .A4(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n659_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n667_), .A3(new_n649_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1325gat));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n313_), .A3(new_n604_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n634_), .A2(new_n501_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(new_n639_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n307_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n634_), .B2(new_n639_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT42), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT42), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1327gat));
  INV_X1    g489(.A(new_n631_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n383_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n652_), .A2(new_n692_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n693_), .A2(G29gat), .A3(new_n635_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n383_), .B1(KEYINPUT105), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n651_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n653_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n629_), .B(new_n699_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n654_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n607_), .A2(KEYINPUT43), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  INV_X1    g502(.A(new_n701_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n650_), .B2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n702_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT105), .B1(new_n695_), .B2(KEYINPUT104), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n607_), .B2(new_n701_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n650_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n707_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n698_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n576_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G29gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n714_), .B2(new_n576_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n694_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  NOR3_X1   g518(.A1(new_n693_), .A2(G36gat), .A3(new_n599_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n712_), .B1(new_n711_), .B2(new_n698_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n697_), .B(new_n707_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n724_), .B(new_n649_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n724_), .B1(new_n714_), .B2(new_n649_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n722_), .B(new_n723_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n649_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT107), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(G36gat), .A3(new_n727_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n723_), .B1(new_n734_), .B2(new_n722_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1329gat));
  INV_X1    g535(.A(new_n693_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G43gat), .B1(new_n737_), .B2(new_n604_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n501_), .A2(new_n447_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n714_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n737_), .B2(new_n685_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n685_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n714_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n291_), .A2(new_n293_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n361_), .A2(new_n365_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n607_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n383_), .A3(new_n691_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n635_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n383_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(new_n704_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n635_), .A2(G57gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1332gat));
  OAI21_X1  g555(.A(G64gat), .B1(new_n750_), .B2(new_n599_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT48), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n599_), .A2(G64gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT109), .Z(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n754_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n750_), .B2(new_n501_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n501_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n754_), .B2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n750_), .B2(new_n639_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n753_), .A2(new_n434_), .A3(new_n685_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n748_), .A2(new_n383_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n711_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n711_), .A2(KEYINPUT111), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(KEYINPUT112), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n576_), .A2(G85gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT113), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n749_), .A2(new_n692_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT110), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n576_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n783_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n781_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n791_), .B2(new_n787_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(G1336gat));
  AOI21_X1  g592(.A(G92gat), .B1(new_n786_), .B2(new_n649_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n649_), .A2(G92gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n779_), .B2(new_n795_), .ZN(G1337gat));
  AOI21_X1  g595(.A(new_n227_), .B1(new_n775_), .B2(new_n604_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n604_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n785_), .A2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OR3_X1    g600(.A1(new_n797_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n786_), .A2(new_n203_), .A3(new_n685_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n711_), .A2(new_n770_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n685_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n808_), .B2(G106gat), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT52), .B(new_n203_), .C1(new_n807_), .C2(new_n685_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n345_), .A2(new_n338_), .A3(new_n331_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n352_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT118), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n336_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n352_), .A4(new_n815_), .ZN(new_n820_));
  AND4_X1   g619(.A1(new_n356_), .A2(new_n283_), .A3(new_n817_), .A4(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n266_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n202_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n284_), .B1(new_n824_), .B2(KEYINPUT55), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n822_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n288_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n821_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n244_), .B1(new_n252_), .B2(new_n224_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n253_), .B1(new_n831_), .B2(KEYINPUT12), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n269_), .A2(new_n273_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(KEYINPUT69), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n202_), .B1(new_n834_), .B2(new_n274_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n278_), .B1(new_n835_), .B2(new_n826_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n827_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n288_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n813_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n830_), .A3(new_n288_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(KEYINPUT58), .A4(new_n821_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n704_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n838_), .A2(new_n845_), .A3(new_n830_), .A4(new_n288_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n830_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n828_), .A2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n746_), .A2(new_n846_), .A3(new_n283_), .A4(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n817_), .A2(new_n356_), .A3(new_n820_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n290_), .A2(new_n850_), .A3(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT119), .B1(new_n290_), .B2(new_n850_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n631_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n844_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n856_), .B(new_n631_), .C1(new_n849_), .C2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n384_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n745_), .A2(new_n366_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n657_), .B2(new_n859_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n291_), .A2(new_n293_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n701_), .A3(new_n862_), .A4(new_n383_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(KEYINPUT54), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT116), .B(new_n865_), .C1(new_n657_), .C2(new_n859_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n635_), .B1(new_n858_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n599_), .A2(new_n641_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n868_), .A2(KEYINPUT120), .A3(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n746_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n858_), .A2(new_n867_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n576_), .A4(new_n870_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n868_), .A2(new_n880_), .A3(KEYINPUT59), .A4(new_n870_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n366_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n878_), .B1(new_n888_), .B2(new_n877_), .ZN(G1340gat));
  AOI21_X1  g688(.A(new_n745_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n745_), .B2(KEYINPUT60), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(KEYINPUT60), .B2(new_n891_), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n890_), .A2(new_n891_), .B1(new_n875_), .B2(new_n893_), .ZN(G1341gat));
  AOI21_X1  g693(.A(G127gat), .B1(new_n876_), .B2(new_n383_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n886_), .A2(new_n887_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n384_), .A2(KEYINPUT123), .ZN(new_n897_));
  MUX2_X1   g696(.A(KEYINPUT123), .B(new_n897_), .S(G127gat), .Z(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n896_), .B2(new_n898_), .ZN(G1342gat));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n876_), .A2(new_n900_), .A3(new_n631_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n886_), .A2(new_n887_), .A3(new_n701_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n900_), .ZN(G1343gat));
  AND3_X1   g702(.A1(new_n868_), .A2(new_n599_), .A3(new_n642_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n746_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n294_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n383_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n904_), .A2(new_n912_), .A3(new_n631_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n904_), .A2(new_n704_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n912_), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n649_), .A2(new_n635_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n501_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n746_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT124), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n685_), .B1(new_n858_), .B2(new_n867_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n471_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n920_), .A2(new_n746_), .A3(new_n537_), .A4(new_n917_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1348gat));
  AND2_X1   g724(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n920_), .A2(new_n917_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n294_), .ZN(new_n930_));
  MUX2_X1   g729(.A(new_n928_), .B(new_n926_), .S(new_n930_), .Z(G1349gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n383_), .ZN(new_n932_));
  MUX2_X1   g731(.A(new_n464_), .B(G183gat), .S(new_n932_), .Z(G1350gat));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n704_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G190gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n929_), .A2(new_n631_), .A3(new_n532_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1351gat));
  AOI211_X1 g736(.A(new_n602_), .B(new_n916_), .C1(new_n858_), .C2(new_n867_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n746_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n294_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n383_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  AND3_X1   g746(.A1(new_n938_), .A2(G218gat), .A3(new_n704_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n938_), .A2(new_n631_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n949_), .A2(KEYINPUT127), .ZN(new_n950_));
  AOI21_X1  g749(.A(G218gat), .B1(new_n949_), .B2(KEYINPUT127), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n948_), .B1(new_n950_), .B2(new_n951_), .ZN(G1355gat));
endmodule


