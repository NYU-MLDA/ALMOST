//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(G204gat), .ZN(new_n203_));
  OAI211_X1 g002(.A(KEYINPUT21), .B(new_n202_), .C1(new_n203_), .C2(G197gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G204gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n203_), .B2(new_n207_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n204_), .B(new_n206_), .C1(new_n209_), .C2(KEYINPUT21), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT92), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n212_), .A2(new_n213_), .B1(G228gat), .B2(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OR4_X1    g016(.A1(KEYINPUT89), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(G141gat), .ZN(new_n219_));
  INV_X1    g018(.A(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(KEYINPUT89), .B2(KEYINPUT3), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n218_), .A2(new_n222_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT86), .ZN(new_n228_));
  INV_X1    g027(.A(G155gat), .ZN(new_n229_));
  INV_X1    g028(.A(G162gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT90), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n227_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n235_), .A2(new_n236_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT87), .B1(new_n235_), .B2(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n239_), .A3(KEYINPUT1), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n221_), .A2(KEYINPUT85), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(KEYINPUT85), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n242_), .A2(new_n243_), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT88), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(KEYINPUT88), .A3(new_n244_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n233_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n212_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n217_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n216_), .B(new_n212_), .C1(new_n249_), .C2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G22gat), .B(G50gat), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n232_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n247_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n245_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n254_), .B1(new_n260_), .B2(KEYINPUT29), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n256_), .B2(new_n261_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n253_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n261_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n262_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n269_), .A2(new_n264_), .B1(new_n252_), .B2(new_n251_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G113gat), .B(G120gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n260_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n246_), .A2(new_n247_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n274_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n258_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n278_), .A3(KEYINPUT4), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n260_), .A2(new_n282_), .A3(new_n274_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n275_), .A2(new_n278_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n280_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G1gat), .B(G29gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G85gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT0), .B(G57gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n279_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT97), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n290_), .B1(new_n285_), .B2(new_n281_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n279_), .A2(KEYINPUT97), .A3(new_n280_), .A4(new_n283_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT95), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n302_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n303_), .B1(new_n306_), .B2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT96), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n303_), .C1(new_n306_), .C2(new_n300_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n308_), .A2(new_n310_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G183gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT94), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(KEYINPUT94), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n316_), .A2(KEYINPUT82), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n316_), .A2(KEYINPUT82), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n314_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n304_), .A2(new_n332_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n328_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n212_), .B1(new_n318_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n324_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT81), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(KEYINPUT81), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n340_), .A2(new_n322_), .A3(new_n341_), .A4(new_n319_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n335_), .A3(new_n317_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n306_), .B1(new_n331_), .B2(new_n311_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n212_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n338_), .A2(KEYINPUT20), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G92gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT18), .B(G64gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n350_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n343_), .A2(new_n344_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n212_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n318_), .A2(new_n337_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n357_), .B(new_n360_), .C1(new_n361_), .C2(new_n212_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n356_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n351_), .B2(new_n362_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n284_), .A2(new_n286_), .A3(KEYINPUT33), .A4(new_n290_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n293_), .A2(new_n299_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n318_), .A2(new_n212_), .A3(new_n337_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n346_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n350_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n338_), .A2(KEYINPUT20), .A3(new_n347_), .A4(new_n357_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT32), .A3(new_n356_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n351_), .A2(new_n362_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n291_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n290_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n374_), .B(new_n376_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n271_), .B1(new_n368_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT31), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n345_), .B(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n274_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n387_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(new_n388_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n359_), .B(new_n384_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT84), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT98), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n355_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n356_), .A2(KEYINPUT98), .ZN(new_n400_));
  AOI211_X1 g199(.A(new_n399_), .B(new_n400_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT99), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n399_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n400_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n373_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT99), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT27), .A4(new_n363_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n395_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n253_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n269_), .A2(new_n252_), .A3(new_n251_), .A4(new_n264_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n396_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n377_), .A2(new_n378_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n380_), .A2(new_n396_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G29gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G43gat), .B(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT15), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G15gat), .B(G22gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G1gat), .A2(G8gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT14), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n424_), .B2(KEYINPUT14), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n423_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G8gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n422_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n431_), .A3(new_n421_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n421_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G113gat), .B(G141gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G169gat), .B(G197gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n447_), .A3(KEYINPUT80), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT12), .ZN(new_n453_));
  AND2_X1   g252(.A1(G57gat), .A2(G64gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G57gat), .A2(G64gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT11), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G57gat), .ZN(new_n457_));
  INV_X1    g256(.A(G64gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G57gat), .A2(G64gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G78gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n456_), .A2(new_n464_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n464_), .B1(new_n456_), .B2(new_n462_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n456_), .A2(new_n464_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT71), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n453_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  AND3_X1   g273(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT67), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT66), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n484_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(G99gat), .B(G106gat), .C1(new_n485_), .C2(KEYINPUT7), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT68), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n484_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n492_), .B(new_n493_), .C1(new_n494_), .C2(new_n484_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n493_), .B1(new_n494_), .B2(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n480_), .A2(new_n481_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n497_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n480_), .B(new_n481_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT10), .B(G99gat), .Z(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT64), .B(G106gat), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n498_), .A2(new_n513_), .A3(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n504_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n473_), .B1(new_n500_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n483_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n486_), .A2(new_n488_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n484_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n492_), .B1(new_n521_), .B2(new_n493_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT68), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .A3(new_n498_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n466_), .A2(new_n526_), .A3(new_n468_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT69), .B1(new_n470_), .B2(new_n471_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n503_), .A2(new_n497_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n517_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n529_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n500_), .B2(new_n516_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n453_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n533_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n534_), .B(KEYINPUT70), .C1(new_n500_), .C2(new_n516_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT73), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n543_), .A2(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(KEYINPUT74), .B2(KEYINPUT13), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n418_), .A2(new_n452_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n230_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT75), .B(G134gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT36), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n422_), .B1(new_n500_), .B2(new_n516_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n525_), .A2(new_n421_), .A3(new_n530_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n567_), .B(new_n570_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n567_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n566_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n572_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT35), .A3(new_n569_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n565_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT76), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n576_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n561_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(KEYINPUT77), .A3(new_n576_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n566_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n561_), .A3(new_n584_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT78), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n589_), .A2(KEYINPUT78), .A3(new_n561_), .A4(new_n584_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n585_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n432_), .B(new_n595_), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n469_), .A2(new_n472_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G211gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT16), .B(G183gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(KEYINPUT17), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n596_), .B(new_n534_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n602_), .B(KEYINPUT17), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n594_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n560_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G1gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n417_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n607_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n589_), .A2(new_n584_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n560_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n417_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(G1324gat));
  INV_X1    g420(.A(new_n410_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G8gat), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT102), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n625_), .B(G8gat), .C1(new_n619_), .C2(new_n622_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(KEYINPUT39), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n628_), .A3(new_n410_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(KEYINPUT102), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n619_), .B2(new_n396_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT41), .Z(new_n636_));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n396_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n611_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(new_n271_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n619_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n611_), .A2(new_n644_), .A3(new_n271_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n380_), .A2(new_n396_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n416_), .A2(new_n417_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n559_), .A2(new_n452_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n617_), .A2(new_n618_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n649_), .A2(KEYINPUT105), .A3(new_n650_), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n417_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n592_), .A2(new_n593_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n585_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT104), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n594_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n659_), .B1(new_n649_), .B2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n418_), .A2(KEYINPUT43), .A3(new_n662_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n650_), .A2(new_n607_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n658_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n649_), .A2(new_n659_), .A3(new_n594_), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n647_), .A2(new_n648_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n659_), .B2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(KEYINPUT44), .A3(new_n607_), .A4(new_n650_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n613_), .ZN(new_n677_));
  MUX2_X1   g476(.A(new_n657_), .B(new_n677_), .S(G29gat), .Z(G1328gat));
  NAND3_X1  g477(.A1(new_n671_), .A2(new_n675_), .A3(new_n410_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n654_), .A2(new_n681_), .A3(new_n410_), .A4(new_n655_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n683_), .A3(KEYINPUT106), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT46), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(KEYINPUT46), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n680_), .A2(new_n683_), .B1(KEYINPUT106), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1329gat));
  NAND3_X1  g488(.A1(new_n676_), .A2(G43gat), .A3(new_n411_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n656_), .B2(new_n396_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g493(.A1(new_n676_), .A2(G50gat), .A3(new_n271_), .ZN(new_n695_));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n656_), .B2(new_n641_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1331gat));
  INV_X1    g497(.A(new_n452_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n418_), .A2(new_n699_), .A3(new_n558_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n608_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n613_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(new_n457_), .A3(new_n417_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1332gat));
  OAI21_X1  g505(.A(G64gat), .B1(new_n704_), .B2(new_n622_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT48), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n458_), .A3(new_n410_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  NAND4_X1  g509(.A1(new_n700_), .A2(new_n617_), .A3(new_n638_), .A4(new_n618_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G71gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n714_), .A3(G71gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n701_), .A2(G71gat), .A3(new_n396_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n713_), .A2(KEYINPUT49), .A3(new_n715_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n704_), .B2(new_n641_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n641_), .A2(G78gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT110), .Z(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n701_), .B2(new_n727_), .ZN(G1335gat));
  AND2_X1   g527(.A1(new_n700_), .A2(new_n651_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  AOI21_X1  g529(.A(G85gat), .B1(new_n730_), .B2(new_n613_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n558_), .A2(new_n699_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n607_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n674_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT112), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n613_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n731_), .B1(new_n737_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n730_), .B2(new_n410_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n736_), .A2(new_n410_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g540(.A1(new_n730_), .A2(new_n510_), .A3(new_n411_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G99gat), .B1(new_n735_), .B2(new_n396_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g544(.A(new_n271_), .B(new_n734_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT113), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n674_), .A2(new_n748_), .A3(new_n271_), .A4(new_n734_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(G106gat), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT52), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n747_), .A2(new_n749_), .A3(new_n752_), .A4(G106gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n730_), .A2(new_n511_), .A3(new_n271_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n758_), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n410_), .A2(new_n417_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n412_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  INV_X1    g564(.A(new_n618_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n452_), .A2(new_n551_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n533_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n537_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n529_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n517_), .B(new_n531_), .C1(new_n771_), .C2(KEYINPUT12), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n769_), .A3(new_n540_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n550_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n777_), .B(new_n549_), .C1(new_n770_), .C2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n767_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n433_), .A2(new_n437_), .A3(new_n435_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n434_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n444_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n447_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n766_), .B1(new_n779_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n765_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT57), .ZN(new_n788_));
  INV_X1    g587(.A(new_n783_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n552_), .B(new_n789_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n769_), .B1(new_n772_), .B2(new_n540_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n772_), .A2(new_n540_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n550_), .B1(new_n795_), .B2(new_n773_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n777_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n550_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n552_), .A4(new_n789_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n792_), .A2(new_n594_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n784_), .B1(new_n799_), .B2(new_n767_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT115), .B(new_n802_), .C1(new_n803_), .C2(new_n766_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n787_), .A2(new_n788_), .A3(new_n801_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n607_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n662_), .A2(new_n558_), .A3(new_n617_), .A4(new_n452_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n608_), .A2(new_n452_), .A3(new_n558_), .A4(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n764_), .B1(new_n806_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n761_), .B1(new_n815_), .B2(new_n452_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n812_), .B1(new_n805_), .B2(new_n607_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT116), .B(KEYINPUT59), .C1(new_n820_), .C2(new_n764_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n764_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n823_));
  OAI21_X1  g622(.A(new_n802_), .B1(new_n803_), .B2(new_n766_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n801_), .A2(new_n788_), .A3(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(new_n607_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n822_), .B(new_n823_), .C1(new_n826_), .C2(new_n812_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n819_), .A2(G113gat), .A3(new_n821_), .A4(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n816_), .B1(new_n828_), .B2(new_n452_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT118), .B(new_n816_), .C1(new_n828_), .C2(new_n452_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1340gat));
  AND2_X1   g632(.A1(new_n819_), .A2(new_n821_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT119), .A3(new_n559_), .A4(new_n827_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n819_), .A2(new_n559_), .A3(new_n821_), .A4(new_n827_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(G120gat), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n814_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n607_), .A2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT120), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(new_n827_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n815_), .B2(new_n607_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n814_), .B2(new_n766_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n834_), .A2(G134gat), .A3(new_n827_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n594_), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n820_), .A2(new_n415_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n762_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n452_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n219_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n558_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n220_), .ZN(G1345gat));
  AND2_X1   g657(.A1(new_n853_), .A2(new_n762_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n617_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n854_), .B2(new_n607_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n863_), .B(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n859_), .B2(new_n766_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n230_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n859_), .B2(new_n868_), .ZN(G1347gat));
  OR2_X1    g668(.A1(new_n826_), .A2(new_n812_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n622_), .A2(new_n613_), .A3(new_n396_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n699_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT122), .Z(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n271_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n301_), .B1(new_n870_), .B2(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT62), .Z(new_n876_));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n641_), .A3(new_n871_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n699_), .A3(new_n305_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1348gat));
  AOI21_X1  g679(.A(G176gat), .B1(new_n878_), .B2(new_n559_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n820_), .A2(new_n271_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n871_), .A2(G176gat), .A3(new_n559_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  AND2_X1   g683(.A1(new_n326_), .A2(new_n327_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n870_), .A2(new_n641_), .A3(new_n885_), .A4(new_n871_), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n886_), .A2(KEYINPUT123), .A3(new_n607_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n607_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n882_), .A2(new_n617_), .A3(new_n871_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n321_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n878_), .A2(new_n319_), .A3(new_n766_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G190gat), .B1(new_n877_), .B2(new_n662_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1351gat));
  NOR2_X1   g693(.A1(new_n622_), .A2(new_n613_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n853_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n452_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n207_), .ZN(G1352gat));
  INV_X1    g697(.A(new_n896_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n559_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G204gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n900_), .B2(new_n203_), .ZN(G1353gat));
  AOI21_X1  g701(.A(new_n896_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n617_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT124), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n904_), .A2(new_n905_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n905_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n903_), .A2(new_n617_), .A3(new_n910_), .A4(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1354gat));
  AOI21_X1  g712(.A(KEYINPUT126), .B1(new_n899_), .B2(new_n766_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT127), .B(G218gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n899_), .A2(KEYINPUT126), .A3(new_n766_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n896_), .A2(new_n662_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n916_), .A2(new_n917_), .B1(new_n915_), .B2(new_n918_), .ZN(G1355gat));
endmodule


