//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT25), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT81), .B1(new_n209_), .B2(G183gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(G183gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT81), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n207_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI211_X1 g017(.A(KEYINPUT82), .B(new_n207_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n221_));
  AND2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT84), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT83), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  INV_X1    g028(.A(new_n222_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n226_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n223_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .A4(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n204_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(KEYINPUT85), .A3(new_n204_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(new_n227_), .A3(new_n222_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n226_), .B2(new_n222_), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n212_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n245_), .A3(new_n206_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n234_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G197gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT93), .B1(new_n248_), .B2(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT93), .ZN(new_n250_));
  INV_X1    g049(.A(G204gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(G197gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(G204gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n253_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(KEYINPUT21), .B2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n257_), .A2(KEYINPUT21), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n256_), .A2(new_n260_), .B1(new_n261_), .B2(new_n254_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n202_), .B1(new_n247_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n222_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n232_), .B1(new_n265_), .B2(new_n229_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n221_), .A2(KEYINPUT84), .A3(new_n222_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n244_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT98), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT98), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n233_), .A2(new_n270_), .A3(new_n244_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n236_), .A2(new_n272_), .A3(new_n206_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n236_), .B2(new_n206_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n208_), .B(KEYINPUT96), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n209_), .A2(G183gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(new_n242_), .A3(new_n207_), .A4(new_n220_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n262_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n264_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT26), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G190gat), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n210_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n288_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n233_), .B1(new_n295_), .B2(KEYINPUT82), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n219_), .A2(new_n220_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n246_), .B(new_n262_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n298_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT95), .B1(new_n298_), .B2(KEYINPUT20), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n262_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n287_), .B1(new_n302_), .B2(new_n286_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n304_));
  XNOR2_X1  g103(.A(G8gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G64gat), .B(G92gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(new_n287_), .C1(new_n302_), .C2(new_n286_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(KEYINPUT100), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n302_), .A2(new_n286_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT100), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n310_), .A4(new_n287_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n286_), .B1(new_n264_), .B2(new_n283_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n286_), .B2(new_n302_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n311_), .B(KEYINPUT27), .C1(new_n319_), .C2(new_n310_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT105), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(KEYINPUT105), .A3(new_n320_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G127gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(G134gat), .ZN(new_n329_));
  INV_X1    g128(.A(G134gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(G127gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT87), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT88), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  INV_X1    g135(.A(G113gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(G120gat), .ZN(new_n338_));
  INV_X1    g137(.A(G120gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(G113gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n342_), .A3(KEYINPUT89), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n342_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n327_), .A2(new_n335_), .A3(new_n332_), .A4(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n346_), .B2(KEYINPUT89), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT31), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n247_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT86), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n354_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n351_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n354_), .A2(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n360_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n354_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n350_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT1), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .A4(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n373_), .A2(new_n377_), .A3(KEYINPUT1), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n373_), .A2(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n370_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n372_), .B(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n380_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n379_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n390_), .A2(KEYINPUT29), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n390_), .B2(KEYINPUT29), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n263_), .B1(new_n389_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n402_), .A2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n400_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n400_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n399_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n396_), .A2(new_n408_), .A3(new_n411_), .A4(new_n398_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n369_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT4), .B1(new_n390_), .B2(new_n347_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n346_), .A2(KEYINPUT101), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT101), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n344_), .A2(new_n345_), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n389_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT102), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n389_), .A2(new_n419_), .A3(KEYINPUT102), .A4(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n390_), .A2(new_n347_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n418_), .B1(new_n427_), .B2(KEYINPUT4), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT0), .ZN(new_n433_));
  INV_X1    g232(.A(G57gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G85gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n422_), .A2(new_n423_), .B1(new_n390_), .B2(new_n347_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n430_), .B1(new_n438_), .B2(new_n425_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n431_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT104), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n439_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT104), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n437_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n437_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n429_), .B(new_n418_), .C1(new_n427_), .C2(KEYINPUT4), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(new_n439_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n417_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n323_), .A2(new_n324_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT106), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT106), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n323_), .A2(new_n450_), .A3(new_n453_), .A4(new_n324_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n449_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(new_n415_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n443_), .B2(new_n437_), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT33), .B(new_n446_), .C1(new_n447_), .C2(new_n439_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n437_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT103), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT103), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n437_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n461_), .B(new_n463_), .C1(new_n430_), .C2(new_n428_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n458_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n312_), .A2(new_n316_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n467_));
  MUX2_X1   g266(.A(new_n319_), .B(new_n303_), .S(new_n467_), .Z(new_n468_));
  AOI22_X1  g267(.A1(new_n465_), .A2(new_n466_), .B1(new_n449_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n456_), .B1(new_n469_), .B2(new_n415_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n369_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n452_), .A2(new_n454_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G190gat), .B(G218gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G134gat), .B(G162gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT36), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT72), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT35), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT34), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT6), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT10), .B(G99gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G85gat), .B(G92gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n496_));
  OAI221_X1 g295(.A(new_n493_), .B1(new_n494_), .B2(G106gat), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n490_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n488_), .A2(KEYINPUT66), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n486_), .A2(new_n502_), .A3(new_n487_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT6), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(KEYINPUT6), .A3(new_n503_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT7), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT67), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n507_), .B(KEYINPUT7), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n495_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n500_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AOI211_X1 g314(.A(KEYINPUT8), .B(new_n495_), .C1(new_n489_), .C2(new_n510_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n499_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n499_), .B(new_n520_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n523_));
  AOI211_X1 g322(.A(new_n479_), .B(new_n482_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n482_), .A2(new_n479_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n482_), .A2(new_n479_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n522_), .A2(new_n526_), .A3(new_n527_), .A4(new_n523_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n478_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(new_n527_), .A3(new_n523_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n525_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n475_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT71), .Z(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n528_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n530_), .A2(KEYINPUT74), .A3(new_n531_), .A4(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n477_), .B(KEYINPUT73), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n537_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT37), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G1gat), .ZN(new_n548_));
  INV_X1    g347(.A(G8gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n551_));
  INV_X1    g350(.A(G15gat), .ZN(new_n552_));
  INV_X1    g351(.A(G22gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G15gat), .A2(G22gat), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n550_), .A2(new_n551_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n551_), .B2(new_n550_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT78), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n557_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT68), .B(G71gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G78gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT11), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(KEYINPUT11), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n566_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n564_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n212_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G211gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n574_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n574_), .A2(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n547_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n506_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n514_), .B1(new_n587_), .B2(new_n504_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n516_), .B1(KEYINPUT8), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n572_), .B1(new_n589_), .B2(new_n498_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n499_), .B(new_n573_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(KEYINPUT12), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n517_), .A2(new_n593_), .A3(new_n572_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n591_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n596_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT69), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n600_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n251_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT5), .B(G176gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n597_), .A2(new_n603_), .A3(new_n600_), .A4(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(KEYINPUT13), .A3(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(KEYINPUT70), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n562_), .B(new_n520_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(G229gat), .A3(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n562_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n521_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n562_), .A2(new_n520_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT79), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT80), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n632_), .B(new_n633_), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n622_), .A2(new_n629_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n472_), .A2(new_n586_), .A3(new_n620_), .A4(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n548_), .A3(new_n449_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(KEYINPUT38), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT107), .Z(new_n644_));
  AND2_X1   g443(.A1(new_n530_), .A2(new_n537_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n472_), .A2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n616_), .A2(new_n584_), .A3(new_n639_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n548_), .B1(new_n648_), .B2(new_n449_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(KEYINPUT38), .B2(new_n642_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n650_), .ZN(G1324gat));
  AND3_X1   g450(.A1(new_n317_), .A2(KEYINPUT105), .A3(new_n320_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT105), .B1(new_n317_), .B2(new_n320_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n640_), .A2(new_n549_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n646_), .A2(new_n655_), .A3(new_n647_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n657_), .A2(new_n658_), .A3(G8gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n657_), .B2(G8gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT108), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n656_), .B(new_n663_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT40), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  AOI21_X1  g468(.A(new_n552_), .B1(new_n648_), .B2(new_n369_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n640_), .A2(new_n552_), .A3(new_n369_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  NAND3_X1  g472(.A1(new_n640_), .A2(new_n553_), .A3(new_n415_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n648_), .A2(new_n415_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G22gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n678_), .A3(G22gat), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(KEYINPUT42), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT42), .B1(new_n677_), .B2(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n680_), .B2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(new_n645_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n616_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n584_), .A3(new_n638_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n472_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n449_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n472_), .B2(new_n547_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n465_), .A2(new_n466_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n449_), .A2(new_n468_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n415_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n321_), .A2(new_n416_), .A3(new_n449_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n471_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n453_), .B1(new_n654_), .B2(new_n450_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n454_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n540_), .A2(new_n541_), .B1(KEYINPUT37), .B2(new_n545_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n685_), .B1(new_n688_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT44), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(G29gat), .A3(new_n449_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n688_), .A2(new_n699_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n685_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n687_), .B1(new_n702_), .B2(new_n705_), .ZN(G1328gat));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n655_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n700_), .A2(KEYINPUT44), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n686_), .A2(new_n710_), .A3(new_n655_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT111), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n711_), .B(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n709_), .B(new_n714_), .C1(KEYINPUT112), .C2(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  INV_X1    g520(.A(G43gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n471_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n700_), .B2(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n705_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G43gat), .B1(new_n686_), .B2(new_n369_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n721_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT113), .B(new_n727_), .C1(new_n705_), .C2(new_n725_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n720_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n701_), .A2(new_n723_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n732_), .B2(new_n708_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n721_), .A3(new_n728_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(KEYINPUT47), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(new_n736_), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n686_), .B2(new_n415_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n701_), .A2(G50gat), .A3(new_n415_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n705_), .ZN(G1331gat));
  NAND4_X1  g539(.A1(new_n646_), .A2(new_n585_), .A3(new_n620_), .A4(new_n639_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n455_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n472_), .A2(new_n586_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n684_), .A2(new_n638_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n449_), .A2(new_n434_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  OR3_X1    g546(.A1(new_n745_), .A2(G64gat), .A3(new_n654_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n741_), .A2(new_n654_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT114), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n752_), .A3(G64gat), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n751_), .A2(KEYINPUT48), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT48), .B1(new_n751_), .B2(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n754_), .B2(new_n755_), .ZN(G1333gat));
  OR3_X1    g555(.A1(new_n745_), .A2(G71gat), .A3(new_n471_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G71gat), .B1(new_n741_), .B2(new_n471_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1334gat));
  OR3_X1    g560(.A1(new_n745_), .A2(G78gat), .A3(new_n416_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n741_), .A2(new_n416_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G78gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT115), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1335gat));
  AOI211_X1 g570(.A(new_n585_), .B(new_n638_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n696_), .A3(new_n645_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n452_), .A2(new_n454_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n683_), .B1(new_n775_), .B2(new_n693_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n772_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n436_), .A3(new_n449_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n744_), .A2(new_n584_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n688_), .B2(new_n699_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n449_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n783_), .B2(new_n436_), .ZN(G1336gat));
  AOI21_X1  g583(.A(G92gat), .B1(new_n779_), .B2(new_n655_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n655_), .A2(G92gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT117), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n782_), .B2(new_n787_), .ZN(G1337gat));
  NOR2_X1   g587(.A1(new_n471_), .A2(new_n494_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n776_), .A2(new_n777_), .A3(new_n772_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n777_), .B1(new_n776_), .B2(new_n772_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n471_), .B(new_n781_), .C1(new_n688_), .C2(new_n699_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n484_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(KEYINPUT120), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n794_), .B2(KEYINPUT51), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n796_), .B1(new_n794_), .B2(KEYINPUT118), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n792_), .B(new_n803_), .C1(new_n793_), .C2(new_n484_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n801_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n484_), .B1(new_n782_), .B2(new_n369_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n789_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT118), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  AND4_X1   g608(.A1(new_n801_), .A2(new_n809_), .A3(KEYINPUT51), .A4(new_n804_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n805_), .B2(new_n810_), .ZN(G1338gat));
  NAND3_X1  g610(.A1(new_n779_), .A2(new_n485_), .A3(new_n415_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n782_), .A2(new_n415_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G106gat), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT52), .B(new_n485_), .C1(new_n782_), .C2(new_n415_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g617(.A1(new_n597_), .A2(KEYINPUT55), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n597_), .A2(KEYINPUT55), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n819_), .A2(new_n820_), .B1(new_n596_), .B2(new_n595_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n609_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n609_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n638_), .A2(new_n611_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n609_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(KEYINPUT122), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n621_), .A2(new_n628_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n634_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n637_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n612_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n683_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n827_), .A2(new_n830_), .B1(new_n612_), .B2(new_n835_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n645_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n609_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n829_), .A3(KEYINPUT123), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n822_), .A2(KEYINPUT123), .A3(new_n823_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n835_), .A2(new_n611_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n842_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n824_), .A2(new_n849_), .A3(new_n826_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n845_), .A4(new_n846_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n698_), .A3(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n838_), .A2(new_n841_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n584_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n614_), .A2(new_n615_), .A3(new_n639_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n586_), .A2(KEYINPUT121), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n698_), .A2(new_n584_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n856_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n855_), .B1(new_n857_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT121), .B1(new_n586_), .B2(new_n856_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n860_), .A3(new_n858_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(KEYINPUT54), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n416_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n655_), .A2(new_n455_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n369_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT124), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n415_), .B1(new_n854_), .B2(new_n867_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  INV_X1    g673(.A(new_n871_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n872_), .A2(new_n337_), .A3(new_n638_), .A4(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n866_), .B1(new_n853_), .B2(new_n584_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n880_), .A2(KEYINPUT59), .A3(new_n415_), .A4(new_n871_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n879_), .A2(new_n881_), .A3(new_n639_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n877_), .B1(new_n882_), .B2(new_n337_), .ZN(G1340gat));
  AOI21_X1  g682(.A(KEYINPUT60), .B1(new_n616_), .B2(new_n339_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(KEYINPUT60), .B2(new_n339_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n872_), .A2(new_n876_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n620_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n879_), .A2(new_n881_), .A3(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(new_n339_), .ZN(G1341gat));
  NAND4_X1  g688(.A1(new_n872_), .A2(new_n328_), .A3(new_n585_), .A4(new_n876_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n879_), .A2(new_n881_), .A3(new_n584_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n328_), .ZN(G1342gat));
  NAND4_X1  g691(.A1(new_n872_), .A2(new_n330_), .A3(new_n645_), .A4(new_n876_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n879_), .A2(new_n881_), .A3(new_n547_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n330_), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n880_), .A2(new_n369_), .A3(new_n416_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n638_), .A3(new_n870_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n620_), .A3(new_n870_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n585_), .A3(new_n870_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  AND4_X1   g702(.A1(G162gat), .A2(new_n896_), .A3(new_n698_), .A4(new_n870_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n369_), .A2(new_n416_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n868_), .A2(new_n645_), .A3(new_n870_), .A4(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(G162gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(KEYINPUT125), .A3(new_n907_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n904_), .B1(new_n910_), .B2(new_n911_), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n654_), .A2(new_n449_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n369_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n873_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT62), .B(G169gat), .C1(new_n916_), .C2(new_n639_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n880_), .A2(new_n415_), .A3(new_n639_), .A4(new_n914_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n203_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n235_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n920_), .A3(new_n921_), .ZN(G1348gat));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n869_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n873_), .A2(KEYINPUT126), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n887_), .A2(new_n914_), .A3(new_n204_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n873_), .A2(new_n616_), .A3(new_n915_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n927_), .B1(new_n204_), .B2(new_n928_), .ZN(G1349gat));
  NOR3_X1   g728(.A1(new_n916_), .A2(new_n584_), .A3(new_n280_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n924_), .A2(new_n585_), .A3(new_n915_), .A4(new_n925_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n212_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n916_), .B2(new_n547_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n645_), .A2(new_n277_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n916_), .B2(new_n934_), .ZN(G1351gat));
  NAND3_X1  g734(.A1(new_n896_), .A2(new_n638_), .A3(new_n913_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g736(.A1(new_n896_), .A2(new_n620_), .A3(new_n913_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT127), .B(G204gat), .Z(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1353gat));
  XNOR2_X1  g739(.A(KEYINPUT63), .B(G211gat), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n896_), .A2(new_n585_), .A3(new_n913_), .A4(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n896_), .A2(new_n913_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n584_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(G1354gat));
  OAI21_X1  g745(.A(G218gat), .B1(new_n943_), .B2(new_n547_), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n683_), .A2(G218gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n943_), .B2(new_n948_), .ZN(G1355gat));
endmodule


