//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  NAND2_X1  g000(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G120gat), .B(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT5), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G176gat), .B(G204gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n209_), .A2(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(KEYINPUT64), .A3(new_n217_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n215_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n216_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n210_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n212_), .A2(new_n214_), .ZN(new_n237_));
  AOI211_X1 g036(.A(KEYINPUT8), .B(new_n231_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n235_), .A3(new_n234_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n231_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n230_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G71gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G78gat), .ZN(new_n245_));
  INV_X1    g044(.A(G78gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G71gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G64gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(KEYINPUT11), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n249_), .B2(KEYINPUT11), .ZN(new_n252_));
  INV_X1    g051(.A(G64gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G57gat), .ZN(new_n254_));
  INV_X1    g053(.A(G57gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G64gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n254_), .A2(new_n256_), .A3(new_n251_), .A4(KEYINPUT11), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n250_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT11), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT65), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n256_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n261_), .A2(new_n264_), .A3(new_n248_), .A4(new_n257_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n243_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT67), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n212_), .A2(new_n214_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n234_), .A2(new_n235_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n241_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT8), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n240_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n259_), .A2(new_n265_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n230_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n243_), .A2(new_n266_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n243_), .A2(KEYINPUT66), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT12), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n243_), .B(new_n266_), .C1(KEYINPUT66), .C2(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n270_), .A2(new_n280_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n268_), .B1(new_n281_), .B2(new_n278_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n207_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n227_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n237_), .B1(new_n208_), .B2(G106gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT12), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n277_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n285_), .ZN(new_n297_));
  AOI211_X1 g096(.A(KEYINPUT67), .B(new_n269_), .C1(new_n292_), .C2(new_n277_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n279_), .B1(new_n278_), .B2(new_n268_), .ZN(new_n299_));
  OAI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n287_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n207_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n288_), .A2(KEYINPUT68), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n288_), .B2(new_n303_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n202_), .B(new_n203_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n288_), .A2(new_n303_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n310_), .A2(KEYINPUT69), .A3(KEYINPUT13), .A4(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G8gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT71), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT71), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G22gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G1gat), .A2(G8gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT14), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n315_), .A2(new_n320_), .A3(new_n318_), .A4(new_n316_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(G231gat), .A3(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(G231gat), .B2(G233gat), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n277_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(G231gat), .ZN(new_n330_));
  INV_X1    g129(.A(G233gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n266_), .B1(new_n332_), .B2(new_n325_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n293_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G127gat), .B(G155gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G183gat), .B(G211gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(KEYINPUT17), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n277_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n266_), .A3(new_n325_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT66), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT73), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n339_), .A2(KEYINPUT17), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n340_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G134gat), .B(G162gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT36), .Z(new_n355_));
  XNOR2_X1  g154(.A(G29gat), .B(G36gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G43gat), .B(G50gat), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT15), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT35), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G232gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT34), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n361_), .A2(new_n243_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n362_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n292_), .A2(new_n360_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n355_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(new_n243_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n365_), .A2(new_n362_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n367_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n354_), .A2(KEYINPUT36), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n370_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(KEYINPUT70), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT37), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n373_), .A2(KEYINPUT70), .A3(KEYINPUT37), .A4(new_n379_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n351_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n313_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G57gat), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G127gat), .B(G134gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT80), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G113gat), .B(G120gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n393_), .A2(KEYINPUT80), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(KEYINPUT80), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT84), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n403_), .A2(KEYINPUT2), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(KEYINPUT2), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .A4(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n402_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G155gat), .A3(G162gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT83), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(KEYINPUT83), .B2(new_n413_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(KEYINPUT1), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n420_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n401_), .B1(new_n416_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n424_), .A3(new_n423_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n420_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n433_), .A2(new_n415_), .A3(new_n400_), .A4(new_n397_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(KEYINPUT4), .A3(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n415_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n401_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n392_), .B(new_n437_), .C1(new_n442_), .C2(new_n436_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n435_), .A2(new_n436_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n391_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(G1gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT100), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT74), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n360_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n358_), .A2(KEYINPUT74), .A3(new_n359_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(new_n324_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n324_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G229gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n361_), .A2(new_n329_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n458_), .B(KEYINPUT75), .Z(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G169gat), .B(G197gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT79), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT30), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT31), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G227gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT78), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(new_n244_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT25), .B(G183gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT76), .B(G190gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT26), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G183gat), .A2(G190gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT23), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(G169gat), .B2(G176gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G169gat), .A2(G176gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT77), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n488_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n485_), .A2(new_n487_), .A3(new_n494_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n481_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n487_), .B1(new_n498_), .B2(G183gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(G169gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n479_), .B(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n401_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n401_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n475_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n474_), .A3(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G226gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT19), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n497_), .A2(new_n502_), .ZN(new_n517_));
  INV_X1    g316(.A(G197gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(G204gat), .ZN(new_n519_));
  INV_X1    g318(.A(G204gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(G197gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT21), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G211gat), .B(G218gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT87), .B1(new_n518_), .B2(G204gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n520_), .A3(G197gat), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n524_), .B(new_n526_), .C1(G197gat), .C2(new_n520_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n522_), .B(new_n523_), .C1(new_n527_), .C2(KEYINPUT21), .ZN(new_n528_));
  INV_X1    g327(.A(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(KEYINPUT21), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n516_), .B1(new_n517_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n490_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n487_), .B1(KEYINPUT24), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT92), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G190gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n480_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n494_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n494_), .A3(KEYINPUT91), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n487_), .B(new_n543_), .C1(KEYINPUT24), .C2(new_n534_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n536_), .A2(new_n541_), .A3(new_n542_), .A4(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546_));
  OR2_X1    g345(.A1(G183gat), .A2(G190gat), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n487_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n487_), .B2(new_n547_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n501_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n531_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n515_), .B1(new_n533_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n503_), .A2(new_n531_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n532_), .A3(new_n550_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT20), .A4(new_n515_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G8gat), .B(G36gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G64gat), .B(G92gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT32), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n443_), .A2(new_n446_), .B1(new_n558_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n533_), .A2(new_n515_), .A3(new_n552_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n533_), .A2(new_n552_), .A3(KEYINPUT99), .A4(new_n515_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n555_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n573_), .A2(new_n574_), .B1(new_n531_), .B2(new_n503_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n555_), .A2(KEYINPUT98), .A3(new_n572_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n515_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n566_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n565_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n391_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n442_), .A2(new_n436_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n435_), .A2(new_n436_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n391_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n580_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n582_), .B1(new_n446_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT20), .B1(new_n503_), .B2(new_n531_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n532_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n514_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n563_), .A3(new_n556_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n563_), .B1(new_n591_), .B2(new_n556_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n588_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n563_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n592_), .A3(KEYINPUT95), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n579_), .B1(new_n587_), .B2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n602_));
  OAI21_X1  g401(.A(G228gat), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n531_), .B2(KEYINPUT88), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n433_), .B2(new_n415_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n606_), .B2(new_n532_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n431_), .A2(new_n432_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n608_));
  OAI221_X1 g407(.A(new_n531_), .B1(KEYINPUT88), .B2(new_n603_), .C1(new_n608_), .C2(new_n605_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G78gat), .B(G106gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n608_), .A2(new_n605_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n608_), .B2(new_n605_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G22gat), .B(G50gat), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n439_), .B2(KEYINPUT29), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n608_), .A2(new_n605_), .A3(new_n614_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n612_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT89), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n624_), .B(new_n611_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n607_), .A2(new_n609_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT89), .B1(new_n628_), .B2(new_n610_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n627_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(KEYINPUT89), .A3(new_n610_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n618_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n620_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n612_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT90), .B1(new_n636_), .B2(new_n629_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n610_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n612_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n635_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n631_), .A2(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n600_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n640_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n627_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n636_), .A2(KEYINPUT90), .A3(new_n629_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT27), .B1(new_n597_), .B2(new_n592_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n596_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n592_), .A2(KEYINPUT27), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n448_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n512_), .B1(new_n642_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n511_), .A2(new_n447_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n641_), .A3(new_n650_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n450_), .B(new_n470_), .C1(new_n652_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n631_), .A2(new_n637_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n447_), .B1(new_n658_), .B2(new_n643_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n659_), .A2(new_n650_), .B1(new_n600_), .B2(new_n641_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n660_), .B2(new_n512_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n450_), .B1(new_n661_), .B2(new_n470_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n386_), .B(new_n449_), .C1(new_n657_), .C2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT101), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n642_), .A2(new_n651_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n655_), .B1(new_n665_), .B2(new_n511_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT100), .B1(new_n666_), .B2(new_n469_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n385_), .B1(new_n667_), .B2(new_n656_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n449_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n307_), .A2(new_n311_), .A3(new_n470_), .A4(new_n351_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n373_), .A2(new_n379_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n661_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n448_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT38), .B1(new_n664_), .B2(new_n670_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT103), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n664_), .A2(new_n670_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n677_), .A4(new_n671_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n680_), .A2(new_n685_), .ZN(G1324gat));
  INV_X1    g485(.A(new_n650_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n674_), .A2(new_n687_), .A3(new_n661_), .A4(new_n675_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G8gat), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(KEYINPUT39), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n650_), .A2(G8gat), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n386_), .B(new_n697_), .C1(new_n657_), .C2(new_n662_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n668_), .A2(KEYINPUT104), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n691_), .A2(new_n692_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n702_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n696_), .A2(new_n702_), .A3(KEYINPUT40), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1325gat));
  OAI21_X1  g508(.A(G15gat), .B1(new_n676_), .B2(new_n511_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT41), .Z(new_n711_));
  INV_X1    g510(.A(new_n668_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n511_), .A2(G15gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1326gat));
  OAI21_X1  g513(.A(G22gat), .B1(new_n676_), .B2(new_n641_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT42), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n641_), .A2(G22gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT107), .Z(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n712_), .B2(new_n718_), .ZN(G1327gat));
  NOR2_X1   g518(.A1(new_n351_), .A2(new_n675_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n313_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n667_), .B2(new_n656_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G29gat), .B1(new_n722_), .B2(new_n447_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n382_), .A2(new_n383_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n724_), .C1(new_n652_), .C2(new_n655_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n312_), .A2(new_n469_), .A3(new_n351_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  INV_X1    g531(.A(new_n730_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n732_), .B(new_n733_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n447_), .A2(G29gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n723_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n735_), .B2(new_n687_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n650_), .A2(G36gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n722_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n722_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n738_), .B1(new_n740_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n745_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n731_), .A2(new_n734_), .A3(new_n650_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n748_), .B(KEYINPUT46), .C1(new_n749_), .C2(new_n739_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  NOR4_X1   g551(.A1(new_n731_), .A2(new_n734_), .A3(new_n752_), .A4(new_n511_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G43gat), .B1(new_n722_), .B2(new_n512_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT47), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n511_), .A2(new_n752_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n735_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n722_), .B2(new_n646_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n646_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n735_), .B2(new_n762_), .ZN(G1331gat));
  INV_X1    g562(.A(new_n351_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n675_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n312_), .A2(new_n469_), .ZN(new_n766_));
  NOR4_X1   g565(.A1(new_n666_), .A2(new_n764_), .A3(new_n765_), .A4(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(G57gat), .A3(new_n447_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT109), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n666_), .A2(new_n470_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n312_), .A2(new_n384_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT108), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n255_), .B1(new_n773_), .B2(new_n448_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n768_), .A2(KEYINPUT109), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1332gat));
  AOI21_X1  g577(.A(new_n253_), .B1(new_n767_), .B2(new_n687_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT48), .Z(new_n780_));
  INV_X1    g579(.A(new_n773_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n253_), .A3(new_n687_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1333gat));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n244_), .A3(new_n512_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n767_), .A2(new_n512_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G71gat), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT49), .B(new_n244_), .C1(new_n767_), .C2(new_n512_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT111), .ZN(G1334gat));
  AOI21_X1  g589(.A(new_n246_), .B1(new_n767_), .B2(new_n646_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT50), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n246_), .A3(new_n646_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1335gat));
  AND2_X1   g593(.A1(new_n312_), .A2(new_n720_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n661_), .A2(new_n469_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n661_), .A2(KEYINPUT112), .A3(new_n469_), .A4(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n223_), .A3(new_n447_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n766_), .A2(new_n351_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n729_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n447_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n804_), .B2(new_n223_), .ZN(G1336gat));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n224_), .A3(new_n687_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n803_), .A2(new_n687_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n224_), .ZN(G1337gat));
  INV_X1    g607(.A(new_n728_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n727_), .B1(new_n661_), .B2(new_n724_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n512_), .B(new_n802_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G99gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G99gat), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n511_), .A2(new_n208_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n800_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n800_), .A2(KEYINPUT114), .A3(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n815_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n813_), .A2(new_n814_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT114), .B1(new_n800_), .B2(new_n817_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n817_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n819_), .B(new_n827_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n824_), .A2(new_n830_), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n800_), .A2(new_n210_), .A3(new_n646_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n729_), .A2(new_n646_), .A3(new_n802_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(G106gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(G106gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT53), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n832_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1339gat));
  NOR2_X1   g640(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n300_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n278_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n269_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n283_), .A2(new_n285_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(KEYINPUT55), .C1(new_n299_), .C2(new_n298_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n207_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n303_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n469_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n267_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n286_), .A2(KEYINPUT55), .B1(new_n268_), .B2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n300_), .A2(new_n844_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT56), .B(new_n207_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n207_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n854_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n460_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n461_), .A2(new_n865_), .A3(new_n456_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n461_), .B2(new_n456_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n462_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n457_), .A2(new_n462_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n466_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n864_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n310_), .B2(new_n304_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n675_), .B(new_n843_), .C1(new_n863_), .C2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n207_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n862_), .A3(new_n858_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n851_), .A2(new_n853_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n873_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n842_), .B1(new_n880_), .B2(new_n765_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n872_), .A2(new_n852_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT58), .B(new_n882_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n724_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n874_), .A2(new_n881_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n764_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n384_), .A2(new_n307_), .A3(new_n469_), .A4(new_n311_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n893_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n687_), .A2(new_n646_), .A3(new_n448_), .A4(new_n511_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(G113gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n470_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(KEYINPUT119), .A3(KEYINPUT59), .ZN(new_n900_));
  OR2_X1    g699(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n896_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n469_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n904_), .B2(new_n898_), .ZN(G1340gat));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n313_), .B2(KEYINPUT60), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n897_), .B(new_n907_), .C1(KEYINPUT60), .C2(new_n906_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n313_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n906_), .ZN(G1341gat));
  INV_X1    g709(.A(G127gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n897_), .A2(new_n911_), .A3(new_n351_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n764_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1342gat));
  INV_X1    g713(.A(G134gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n897_), .A2(new_n915_), .A3(new_n765_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n725_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1343gat));
  NOR4_X1   g717(.A1(new_n687_), .A2(new_n641_), .A3(new_n512_), .A4(new_n448_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n894_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n470_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n313_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT120), .B(G148gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n764_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  OR3_X1    g728(.A1(new_n920_), .A2(G162gat), .A3(new_n675_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G162gat), .B1(new_n920_), .B2(new_n725_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1347gat));
  INV_X1    g731(.A(KEYINPUT22), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n687_), .A2(new_n653_), .A3(new_n641_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n894_), .A2(new_n933_), .A3(new_n470_), .A4(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(G169gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n936_), .A2(KEYINPUT62), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n892_), .B1(new_n888_), .B2(new_n764_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(new_n469_), .A3(new_n934_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n933_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n894_), .A2(new_n939_), .A3(new_n470_), .A4(new_n935_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G169gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n938_), .B1(new_n942_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(KEYINPUT121), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n947_), .B(new_n938_), .C1(new_n942_), .C2(new_n944_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1348gat));
  NOR2_X1   g748(.A1(new_n940_), .A2(new_n934_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n312_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT122), .B(G176gat), .Z(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1349gat));
  NAND2_X1  g752(.A1(new_n950_), .A2(new_n351_), .ZN(new_n954_));
  MUX2_X1   g753(.A(new_n480_), .B(G183gat), .S(new_n954_), .Z(G1350gat));
  NAND3_X1  g754(.A1(new_n950_), .A2(new_n537_), .A3(new_n765_), .ZN(new_n956_));
  INV_X1    g755(.A(G190gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n940_), .A2(new_n725_), .A3(new_n934_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n956_), .B1(new_n957_), .B2(new_n958_), .ZN(G1351gat));
  NAND3_X1  g758(.A1(new_n659_), .A2(new_n687_), .A3(new_n511_), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n894_), .A2(new_n470_), .A3(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(KEYINPUT124), .B1(new_n962_), .B2(new_n518_), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT123), .B1(new_n962_), .B2(new_n518_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n940_), .A2(new_n960_), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966_));
  NAND4_X1  g765(.A1(new_n965_), .A2(new_n966_), .A3(G197gat), .A4(new_n470_), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n963_), .A2(new_n964_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n964_), .B1(new_n963_), .B2(new_n967_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n965_), .A2(new_n312_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g771(.A1(new_n940_), .A2(new_n764_), .A3(new_n960_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974_));
  OR2_X1    g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  OR3_X1    g774(.A1(new_n973_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n974_), .B1(new_n973_), .B2(new_n975_), .ZN(new_n977_));
  XOR2_X1   g776(.A(KEYINPUT63), .B(G211gat), .Z(new_n978_));
  AOI22_X1  g777(.A1(new_n976_), .A2(new_n977_), .B1(new_n973_), .B2(new_n978_), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n965_), .B2(new_n765_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n724_), .A2(G218gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(KEYINPUT126), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n980_), .B1(new_n965_), .B2(new_n982_), .ZN(G1355gat));
endmodule


