//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  AOI22_X1  g007(.A1(new_n203_), .A2(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n213_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n210_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n221_), .A2(KEYINPUT64), .A3(new_n217_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n209_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n206_), .A2(new_n208_), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n206_), .A2(new_n208_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n214_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT65), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n224_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT65), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n224_), .B1(new_n241_), .B2(new_n236_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n233_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n225_), .A2(new_n231_), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n223_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G64gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n249_));
  XOR2_X1   g048(.A(G71gat), .B(G78gat), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n223_), .B(new_n253_), .C1(new_n240_), .C2(new_n245_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n257_), .B(new_n258_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n259_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G230gat), .A3(G233gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT5), .B(G176gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT69), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n267_), .A2(new_n272_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n267_), .A2(KEYINPUT69), .A3(new_n272_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT74), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G43gat), .B(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n294_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n283_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n294_), .B(new_n297_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT78), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n294_), .A2(new_n297_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n297_), .B(KEYINPUT15), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n300_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT79), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n305_), .A2(new_n310_), .A3(new_n300_), .A4(new_n307_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n301_), .A2(new_n304_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G169gat), .B(G197gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n282_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G227gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(G71gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G15gat), .B(G43gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT22), .B(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(G176gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(G183gat), .C2(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G190gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT80), .B1(new_n347_), .B2(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350_));
  INV_X1    g149(.A(G190gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT26), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n346_), .A2(new_n348_), .A3(new_n349_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT81), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n349_), .A2(new_n352_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n336_), .A2(new_n337_), .ZN(new_n359_));
  OR3_X1    g158(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n339_), .B(KEYINPUT82), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n359_), .B(new_n360_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n343_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT30), .B1(new_n368_), .B2(new_n343_), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n330_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n365_), .A2(new_n366_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n368_), .A2(KEYINPUT30), .A3(new_n343_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n370_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n329_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT85), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n374_), .A2(new_n379_), .A3(new_n380_), .A4(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n374_), .A2(new_n380_), .A3(new_n379_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n385_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n380_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n386_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  INV_X1    g192(.A(G141gat), .ZN(new_n394_));
  INV_X1    g193(.A(G148gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT87), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(KEYINPUT1), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(KEYINPUT1), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT88), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n393_), .B(new_n396_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(KEYINPUT3), .ZN(new_n404_));
  OR3_X1    g203(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(KEYINPUT2), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n404_), .B(new_n405_), .C1(new_n393_), .C2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(KEYINPUT2), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n409_), .A2(new_n410_), .B1(G141gat), .B2(G148gat), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n398_), .B(new_n399_), .C1(new_n408_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n403_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(KEYINPUT29), .ZN(new_n414_));
  XOR2_X1   g213(.A(G78gat), .B(G106gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G211gat), .B(G218gat), .Z(new_n418_));
  OAI21_X1  g217(.A(new_n269_), .B1(KEYINPUT91), .B2(G197gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT90), .B(G204gat), .ZN(new_n420_));
  INV_X1    g219(.A(G197gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(KEYINPUT91), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n423_), .B2(KEYINPUT21), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(G197gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(G204gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n426_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n418_), .A2(KEYINPUT21), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n424_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n413_), .B2(KEYINPUT29), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT28), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n432_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n417_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n416_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n392_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n383_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n382_), .B(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n403_), .A3(new_n412_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n413_), .A2(new_n384_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT4), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n413_), .A2(new_n384_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT99), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(new_n213_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT0), .B(G57gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n446_), .A2(new_n447_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n449_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n448_), .A2(new_n460_), .A3(new_n451_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT98), .A4(new_n449_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n463_), .A2(new_n466_), .A3(new_n458_), .A4(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n424_), .A2(new_n428_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n430_), .A2(new_n429_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n351_), .A2(KEYINPUT26), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n348_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT92), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n348_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n478_), .A2(new_n480_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n339_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n359_), .B(new_n360_), .C1(new_n482_), .C2(new_n362_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n342_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT20), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n475_), .B(KEYINPUT95), .C1(new_n343_), .C2(new_n368_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n365_), .B2(new_n431_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n485_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT19), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n489_), .A2(KEYINPUT96), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT96), .B1(new_n489_), .B2(new_n492_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495_));
  INV_X1    g294(.A(new_n484_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n431_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n475_), .A2(KEYINPUT93), .A3(new_n484_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n365_), .A2(new_n431_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n497_), .A2(KEYINPUT20), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n500_), .A2(KEYINPUT94), .A3(new_n491_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT94), .B1(new_n500_), .B2(new_n491_), .ZN(new_n502_));
  OAI22_X1  g301(.A1(new_n493_), .A2(new_n494_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G8gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n211_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT18), .B(G64gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n489_), .A2(new_n492_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n489_), .A2(KEYINPUT96), .A3(new_n492_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n500_), .A2(new_n491_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n500_), .A2(KEYINPUT94), .A3(new_n491_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n508_), .A2(new_n520_), .A3(KEYINPUT97), .ZN(new_n521_));
  OR3_X1    g320(.A1(new_n503_), .A2(KEYINPUT97), .A3(new_n507_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n472_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n463_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n457_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n468_), .ZN(new_n527_));
  OR3_X1    g326(.A1(new_n524_), .A2(new_n526_), .A3(new_n457_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n503_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n500_), .A2(new_n491_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n492_), .B2(new_n489_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(new_n530_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n529_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n443_), .B1(new_n523_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n521_), .A2(new_n522_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n391_), .A2(new_n442_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n441_), .B(new_n386_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n533_), .B2(new_n507_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n520_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n541_), .A3(new_n529_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n322_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G127gat), .B(G155gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G211gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n292_), .A2(new_n293_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n253_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n293_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n289_), .A2(new_n291_), .ZN(new_n555_));
  OAI211_X1 g354(.A(G231gat), .B(G233gat), .C1(new_n554_), .C2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n292_), .A2(new_n293_), .A3(new_n550_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n254_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n549_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  AOI211_X1 g361(.A(G211gat), .B(new_n562_), .C1(new_n553_), .C2(new_n558_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n548_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n551_), .A2(new_n552_), .A3(new_n253_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n254_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n560_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G211gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n549_), .A3(new_n560_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n547_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT16), .B(G183gat), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n573_));
  NAND3_X1  g372(.A1(new_n553_), .A2(new_n558_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT77), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT77), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n574_), .A4(new_n572_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n246_), .A2(new_n306_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n582_), .B(new_n585_), .C1(new_n298_), .C2(new_n246_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT70), .Z(new_n588_));
  AND2_X1   g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n586_), .A2(new_n588_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT71), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT36), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n589_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n594_), .ZN(new_n597_));
  OAI22_X1  g396(.A1(new_n589_), .A2(new_n590_), .B1(KEYINPUT36), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT101), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n546_), .A2(new_n581_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n529_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n202_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT72), .B1(new_n596_), .B2(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n577_), .A2(new_n580_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n546_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n202_), .A3(new_n605_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT103), .B1(new_n618_), .B2(new_n606_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1324gat));
  NAND2_X1  g419(.A1(new_n538_), .A2(new_n543_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n613_), .A2(new_n284_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT104), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n602_), .A2(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G8gat), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT40), .B(new_n623_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  NAND2_X1  g431(.A1(new_n604_), .A2(new_n392_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G15gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n636_), .A3(G15gat), .ZN(new_n637_));
  NOR4_X1   g436(.A1(new_n546_), .A2(G15gat), .A3(new_n391_), .A4(new_n612_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT105), .Z(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n637_), .A3(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n613_), .A2(new_n641_), .A3(new_n442_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n604_), .A2(new_n442_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(G22gat), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT42), .B(new_n641_), .C1(new_n604_), .C2(new_n442_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  XNOR2_X1  g446(.A(new_n608_), .B(KEYINPUT37), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n545_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT43), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n545_), .A2(new_n651_), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n581_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n282_), .A3(new_n321_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(KEYINPUT44), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n605_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G29gat), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n322_), .A2(new_n545_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n654_), .A2(new_n600_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n529_), .A2(G29gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT106), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n663_), .B2(new_n665_), .ZN(G1328gat));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n621_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G36gat), .B1(new_n657_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n621_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n661_), .A2(new_n662_), .A3(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT45), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT107), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(KEYINPUT107), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n668_), .A2(KEYINPUT107), .A3(new_n674_), .A4(new_n672_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  INV_X1    g478(.A(G43gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n663_), .B2(new_n391_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n658_), .A2(G43gat), .A3(new_n392_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n657_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT47), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n683_), .B(new_n687_), .C1(new_n657_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1330gat));
  INV_X1    g488(.A(new_n663_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G50gat), .B1(new_n690_), .B2(new_n442_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n657_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n658_), .A2(G50gat), .A3(new_n442_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(G1331gat));
  AOI21_X1  g493(.A(new_n320_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n282_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(new_n654_), .A3(new_n600_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(G57gat), .A3(new_n605_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n282_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n612_), .A2(new_n700_), .A3(KEYINPUT109), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT109), .B1(new_n612_), .B2(new_n700_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n695_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n704_), .B2(new_n529_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n705_), .B2(KEYINPUT110), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(KEYINPUT110), .B2(new_n705_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n697_), .B2(new_n621_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT48), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n708_), .A3(new_n621_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1333gat));
  AOI21_X1  g511(.A(new_n324_), .B1(new_n697_), .B2(new_n392_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT49), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n703_), .A2(new_n324_), .A3(new_n392_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n697_), .B2(new_n442_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT50), .Z(new_n719_));
  NAND2_X1  g518(.A1(new_n442_), .A2(new_n717_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT111), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n704_), .B2(new_n721_), .ZN(G1335gat));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n650_), .A2(new_n723_), .A3(new_n652_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n651_), .B1(new_n545_), .B2(new_n648_), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT43), .B(new_n610_), .C1(new_n536_), .C2(new_n544_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT112), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n282_), .A2(new_n321_), .A3(new_n581_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n732_), .B(new_n729_), .C1(new_n724_), .C2(new_n727_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n529_), .A2(new_n213_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n696_), .A2(new_n605_), .A3(new_n662_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n734_), .A2(new_n735_), .B1(new_n213_), .B2(new_n736_), .ZN(G1336gat));
  NAND3_X1  g536(.A1(new_n696_), .A2(new_n621_), .A3(new_n662_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n211_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT114), .Z(new_n740_));
  NOR2_X1   g539(.A1(new_n669_), .A2(new_n211_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n734_), .B2(new_n741_), .ZN(G1337gat));
  NAND2_X1  g541(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n326_), .B1(new_n734_), .B2(new_n392_), .ZN(new_n745_));
  AND4_X1   g544(.A1(new_n203_), .A2(new_n696_), .A3(new_n392_), .A4(new_n662_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT115), .Z(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n731_), .A2(new_n733_), .A3(new_n391_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n749_), .B(new_n743_), .C1(new_n750_), .C2(new_n326_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1338gat));
  NAND4_X1  g551(.A1(new_n696_), .A2(new_n204_), .A3(new_n442_), .A4(new_n662_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n653_), .A2(new_n442_), .A3(new_n730_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G106gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  INV_X1    g559(.A(new_n319_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n318_), .B1(new_n302_), .B2(new_n300_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n305_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR4_X1   g563(.A1(new_n276_), .A2(new_n761_), .A3(new_n277_), .A4(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n272_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT118), .B1(new_n264_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n259_), .A2(new_n261_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT68), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n246_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT12), .B1(new_n246_), .B2(new_n254_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n772_), .A2(new_n775_), .A3(new_n776_), .A4(KEYINPUT55), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n264_), .A2(new_n778_), .A3(new_n767_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n768_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n257_), .A2(new_n258_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n259_), .ZN(new_n782_));
  OAI211_X1 g581(.A(G230gat), .B(G233gat), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT55), .B1(new_n772_), .B2(new_n775_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n778_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n766_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT120), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n787_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT56), .B(new_n766_), .C1(new_n780_), .C2(new_n785_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n320_), .A2(new_n273_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n765_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n760_), .B1(new_n796_), .B2(new_n601_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n768_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n785_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n272_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n788_), .A2(KEYINPUT120), .B1(new_n800_), .B2(KEYINPUT56), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n794_), .B1(new_n801_), .B2(new_n791_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT57), .B(new_n600_), .C1(new_n802_), .C2(new_n765_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n764_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n273_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n786_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n807_), .B2(new_n792_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n648_), .B1(new_n808_), .B2(KEYINPUT58), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n810_), .B(new_n805_), .C1(new_n807_), .C2(new_n792_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n797_), .A2(new_n803_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n581_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n320_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n611_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n611_), .B2(new_n817_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n540_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n621_), .A2(new_n529_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n320_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n828_), .A3(new_n823_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n320_), .A2(G113gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(G1340gat));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n700_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n825_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n827_), .A2(new_n282_), .A3(new_n829_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g636(.A(G127gat), .B1(new_n825_), .B2(new_n654_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n654_), .A2(G127gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n830_), .B2(new_n839_), .ZN(G1342gat));
  AOI21_X1  g639(.A(G134gat), .B1(new_n825_), .B2(new_n601_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n648_), .A2(G134gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT121), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n830_), .B2(new_n843_), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n820_), .B1(new_n581_), .B2(new_n814_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n539_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n823_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n321_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n394_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n700_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n395_), .ZN(G1345gat));
  NOR2_X1   g650(.A1(new_n847_), .A2(new_n581_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n852_), .B(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(new_n847_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G162gat), .B1(new_n856_), .B2(new_n601_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n648_), .A2(G162gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT122), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n856_), .B2(new_n859_), .ZN(G1347gat));
  XOR2_X1   g659(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n861_));
  INV_X1    g660(.A(new_n540_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n669_), .A2(new_n605_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n600_), .B1(new_n802_), .B2(new_n765_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n812_), .B1(new_n864_), .B2(new_n760_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n654_), .B1(new_n865_), .B2(new_n803_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n862_), .B(new_n863_), .C1(new_n866_), .C2(new_n820_), .ZN(new_n867_));
  OAI211_X1 g666(.A(G169gat), .B(new_n861_), .C1(new_n867_), .C2(new_n321_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n822_), .A2(new_n320_), .A3(new_n331_), .A4(new_n863_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n822_), .A2(new_n320_), .A3(new_n863_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n861_), .B1(new_n871_), .B2(G169gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT124), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n861_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n863_), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n845_), .A2(new_n321_), .A3(new_n540_), .A4(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G169gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n874_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n869_), .A4(new_n868_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n873_), .A2(new_n880_), .ZN(G1348gat));
  XNOR2_X1  g680(.A(KEYINPUT125), .B(G176gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n332_), .A2(KEYINPUT125), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n867_), .A2(new_n700_), .ZN(new_n884_));
  MUX2_X1   g683(.A(new_n882_), .B(new_n883_), .S(new_n884_), .Z(G1349gat));
  NOR2_X1   g684(.A1(new_n867_), .A2(new_n581_), .ZN(new_n886_));
  MUX2_X1   g685(.A(G183gat), .B(new_n346_), .S(new_n886_), .Z(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n867_), .B2(new_n610_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n478_), .A2(new_n480_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n601_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n867_), .B2(new_n890_), .ZN(G1351gat));
  NOR3_X1   g690(.A1(new_n845_), .A2(new_n539_), .A3(new_n875_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n320_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n282_), .ZN(new_n895_));
  MUX2_X1   g694(.A(new_n420_), .B(G204gat), .S(new_n895_), .Z(G1353gat));
  AOI211_X1 g695(.A(KEYINPUT63), .B(G211gat), .C1(new_n892_), .C2(new_n654_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n892_), .A2(new_n654_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT63), .B(G211gat), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1354gat));
  XOR2_X1   g699(.A(KEYINPUT126), .B(G218gat), .Z(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n648_), .A3(new_n901_), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n845_), .A2(new_n539_), .A3(new_n600_), .A4(new_n875_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n901_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n902_), .B(new_n906_), .C1(new_n903_), .C2(new_n901_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1355gat));
endmodule


