//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  NOR2_X1   g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT89), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n202_), .B1(new_n207_), .B2(G204gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n204_), .A2(new_n206_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n209_), .B1(new_n208_), .B2(KEYINPUT21), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n212_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT92), .ZN(new_n222_));
  INV_X1    g021(.A(new_n202_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT89), .B(G197gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n213_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n210_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n209_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n212_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G155gat), .B(G162gat), .Z(new_n230_));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT86), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234_));
  INV_X1    g033(.A(G141gat), .ZN(new_n235_));
  INV_X1    g034(.A(G148gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n231_), .B2(KEYINPUT86), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n230_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT87), .B(new_n230_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n235_), .A2(new_n236_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n231_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n230_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n222_), .A2(new_n229_), .B1(new_n252_), .B2(KEYINPUT29), .ZN(new_n253_));
  INV_X1    g052(.A(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT88), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G228gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(G228gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT93), .B1(new_n253_), .B2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n227_), .A2(new_n228_), .A3(new_n212_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n228_), .B1(new_n227_), .B2(new_n212_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n250_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n262_), .A2(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT93), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n259_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n221_), .A2(new_n260_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n259_), .B1(new_n227_), .B2(new_n212_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(KEYINPUT91), .C1(new_n264_), .C2(new_n265_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G78gat), .B(G106gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n261_), .A2(new_n268_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT94), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n265_), .A2(new_n264_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G22gat), .B(G50gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT28), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n280_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n261_), .A2(new_n268_), .A3(new_n275_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n276_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n278_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT95), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(new_n290_), .A3(new_n283_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G226gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT19), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT20), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n262_), .A2(new_n263_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT22), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G169gat), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT22), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT99), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT99), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n313_), .A3(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n314_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT96), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n320_), .A2(KEYINPUT26), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(KEYINPUT26), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT96), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT25), .B(G183gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT81), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G169gat), .B2(G176gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n333_), .A2(new_n335_), .A3(KEYINPUT24), .A4(new_n310_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(KEYINPUT97), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n332_), .A2(KEYINPUT81), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n334_), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT98), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n317_), .A2(new_n318_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT24), .B1(new_n333_), .B2(new_n335_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT98), .B1(new_n346_), .B2(new_n343_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT97), .B1(new_n331_), .B2(new_n336_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n323_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n301_), .B1(new_n302_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT103), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n330_), .A2(new_n328_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n341_), .A2(new_n354_), .A3(new_n336_), .A4(new_n344_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n306_), .A2(KEYINPUT82), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n306_), .A2(KEYINPUT82), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n308_), .A4(new_n304_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n310_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n355_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n352_), .A2(new_n353_), .B1(new_n221_), .B2(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n350_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT103), .B1(new_n364_), .B2(new_n301_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n300_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n218_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n209_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n225_), .B2(new_n210_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n369_), .A2(new_n371_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n331_), .A2(new_n336_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n345_), .A2(new_n347_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n337_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n377_), .B2(new_n323_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n221_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n378_), .A2(new_n299_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n297_), .B1(new_n366_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n372_), .A3(new_n323_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n301_), .B1(new_n362_), .B2(new_n221_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n300_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n350_), .A2(new_n221_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n379_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n299_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n382_), .B1(new_n390_), .B2(new_n296_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n378_), .A2(new_n300_), .A3(new_n379_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n299_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n296_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n386_), .A2(new_n389_), .A3(new_n297_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n382_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT104), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT104), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n399_), .A3(new_n382_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n381_), .A2(new_n391_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n362_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G43gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G15gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n408_), .B(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT84), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n402_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G134gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G127gat), .ZN(new_n418_));
  INV_X1    g217(.A(G127gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G134gat), .ZN(new_n420_));
  INV_X1    g219(.A(G120gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G113gat), .ZN(new_n422_));
  INV_X1    g221(.A(G113gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G120gat), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n418_), .A2(new_n420_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n418_), .A2(new_n420_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT31), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n412_), .A2(new_n402_), .A3(new_n415_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n428_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n432_), .B2(new_n416_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n252_), .A2(new_n427_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n265_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(KEYINPUT4), .A3(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n265_), .A2(KEYINPUT4), .A3(new_n440_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n438_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n437_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n265_), .A2(new_n440_), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n427_), .B(new_n250_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n446_), .B1(new_n452_), .B2(new_n443_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n437_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n448_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n433_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n290_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n283_), .ZN(new_n460_));
  AOI211_X1 g259(.A(KEYINPUT95), .B(new_n460_), .C1(new_n278_), .C2(KEYINPUT94), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n288_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  AND4_X1   g261(.A1(new_n292_), .A2(new_n401_), .A3(new_n458_), .A4(new_n462_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n449_), .A2(new_n450_), .A3(new_n438_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT101), .B1(new_n464_), .B2(new_n437_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n442_), .A2(new_n438_), .A3(new_n444_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n439_), .A2(new_n446_), .A3(new_n441_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT101), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n454_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n470_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT33), .B1(new_n472_), .B2(KEYINPUT100), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n448_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n471_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT102), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT102), .A4(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n390_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n352_), .A2(new_n353_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n362_), .A2(new_n221_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n365_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n380_), .B1(new_n485_), .B2(new_n299_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n457_), .B(new_n482_), .C1(new_n486_), .C2(new_n481_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n480_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n292_), .A3(new_n462_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n292_), .A2(new_n462_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n457_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n401_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n463_), .B1(new_n493_), .B2(new_n433_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT10), .B(G99gat), .Z(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G85gat), .B(G92gat), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT9), .ZN(new_n500_));
  INV_X1    g299(.A(G85gat), .ZN(new_n501_));
  INV_X1    g300(.A(G92gat), .ZN(new_n502_));
  OR3_X1    g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT9), .ZN(new_n503_));
  INV_X1    g302(.A(G99gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT6), .B1(new_n504_), .B2(new_n497_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n498_), .A2(new_n500_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT65), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  NOR2_X1   g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(KEYINPUT64), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT64), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n514_), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(KEYINPUT64), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT65), .A4(new_n511_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n504_), .A2(new_n497_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n505_), .A2(new_n507_), .B1(new_n520_), .B2(KEYINPUT7), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n499_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n522_), .B2(new_n499_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n509_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n495_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n532_));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n522_), .A2(new_n499_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT8), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n522_), .A2(new_n523_), .A3(new_n499_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n536_), .B1(new_n540_), .B2(new_n509_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n509_), .B(new_n536_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n528_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n509_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT12), .B1(new_n546_), .B2(KEYINPUT66), .ZN(new_n547_));
  INV_X1    g346(.A(new_n536_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n526_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n544_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(G230gat), .B(G233gat), .C1(new_n541_), .C2(new_n543_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT68), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G176gat), .B(G204gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n552_), .A2(new_n553_), .A3(new_n560_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT69), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n554_), .A2(new_n565_), .A3(new_n561_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT74), .B(G15gat), .ZN(new_n572_));
  INV_X1    g371(.A(G22gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G1gat), .ZN(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G1gat), .B(G8gat), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n579_), .A3(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G43gat), .B(G50gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G29gat), .B(G36gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n587_), .B(KEYINPUT15), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n583_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n589_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n587_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n593_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n594_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n583_), .A2(new_n587_), .ZN(new_n602_));
  OAI211_X1 g401(.A(G229gat), .B(G233gat), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n589_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n598_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT79), .B1(new_n600_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n599_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT79), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n494_), .A2(new_n571_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n590_), .A2(new_n526_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT71), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT34), .Z(new_n618_));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n615_), .B(new_n620_), .C1(new_n526_), .C2(new_n587_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n619_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G190gat), .B(G218gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT70), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT36), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT72), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n623_), .A2(new_n630_), .A3(new_n624_), .A4(new_n629_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(KEYINPUT37), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT73), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n632_), .A3(KEYINPUT73), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n634_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n583_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n583_), .A2(new_n644_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n536_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n583_), .A2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n583_), .A2(new_n644_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n548_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n527_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n536_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n548_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(KEYINPUT66), .ZN(new_n654_));
  XOR2_X1   g453(.A(G127gat), .B(G155gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(G183gat), .B(G211gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT17), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT76), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n651_), .A2(new_n654_), .A3(new_n661_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n659_), .A2(KEYINPUT17), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n652_), .A2(new_n653_), .A3(new_n660_), .A4(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(KEYINPUT77), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT77), .B1(new_n662_), .B2(new_n664_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT78), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n667_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT78), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n665_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n643_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n614_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n575_), .A3(new_n457_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT38), .ZN(new_n677_));
  INV_X1    g476(.A(new_n640_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n494_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n666_), .A2(new_n667_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n611_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n571_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G1gat), .B1(new_n683_), .B2(new_n491_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n677_), .A2(new_n684_), .ZN(G1324gat));
  OAI21_X1  g484(.A(G8gat), .B1(new_n683_), .B2(new_n401_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(new_n401_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n675_), .A2(new_n576_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n683_), .B2(new_n433_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n433_), .A2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n674_), .B2(new_n696_), .ZN(G1326gat));
  INV_X1    g496(.A(new_n490_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G22gat), .B1(new_n683_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n675_), .A2(new_n573_), .A3(new_n490_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1327gat));
  INV_X1    g501(.A(new_n672_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n640_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n614_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n457_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n494_), .B2(new_n642_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n433_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT107), .B(new_n643_), .C1(new_n711_), .C2(new_n463_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(KEYINPUT43), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n708_), .B(new_n714_), .C1(new_n494_), .C2(new_n642_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n713_), .A2(new_n672_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n682_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n457_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n707_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n688_), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n705_), .A2(G36gat), .A3(new_n401_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT45), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(KEYINPUT46), .A3(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  NAND4_X1  g531(.A1(new_n719_), .A2(G43gat), .A3(new_n710_), .A4(new_n720_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n705_), .A2(new_n433_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(G43gat), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n706_), .B2(new_n490_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n490_), .A2(G50gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n721_), .B2(new_n738_), .ZN(G1331gat));
  NAND3_X1  g538(.A1(new_n613_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n679_), .A2(new_n571_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n491_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n494_), .A2(new_n570_), .A3(new_n611_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n673_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n491_), .A2(G57gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  OAI21_X1  g546(.A(G64gat), .B1(new_n742_), .B2(new_n401_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  NOR3_X1   g548(.A1(new_n745_), .A2(G64gat), .A3(new_n401_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT108), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n742_), .B2(new_n433_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n433_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n745_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n742_), .B2(new_n698_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n698_), .A2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n745_), .B2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n744_), .A2(new_n704_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n501_), .A3(new_n457_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n570_), .A2(new_n611_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n713_), .A2(new_n672_), .A3(new_n715_), .A4(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n715_), .A2(new_n672_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(KEYINPUT109), .A3(new_n713_), .A4(new_n764_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(KEYINPUT110), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT110), .B1(new_n767_), .B2(new_n769_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n491_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n763_), .B1(new_n772_), .B2(new_n501_), .ZN(G1336gat));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n502_), .A3(new_n688_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n770_), .A2(new_n771_), .A3(new_n401_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n502_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT111), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n774_), .C1(new_n775_), .C2(new_n502_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1337gat));
  AOI21_X1  g579(.A(new_n433_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n710_), .A2(new_n496_), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n781_), .A2(new_n504_), .B1(new_n761_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g583(.A1(new_n762_), .A2(new_n497_), .A3(new_n490_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n786_));
  NOR2_X1   g585(.A1(new_n765_), .A2(new_n698_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n497_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT112), .B1(new_n765_), .B2(new_n698_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n716_), .A2(new_n788_), .A3(new_n490_), .A4(new_n764_), .ZN(new_n792_));
  AND4_X1   g591(.A1(G106gat), .A2(new_n792_), .A3(new_n790_), .A4(new_n786_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n785_), .B(new_n795_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n643_), .A2(new_n740_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n570_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(new_n570_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n592_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n589_), .A2(new_n591_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n805_), .B(new_n599_), .C1(new_n592_), .C2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n608_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n564_), .A2(KEYINPUT115), .A3(new_n566_), .A4(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n564_), .A2(new_n566_), .A3(new_n808_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n551_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n552_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n544_), .A2(new_n550_), .A3(KEYINPUT55), .A4(new_n551_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n561_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n560_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n611_), .A2(new_n563_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n809_), .B(new_n812_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n640_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n817_), .A2(new_n561_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n819_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n808_), .A2(new_n563_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n818_), .B2(KEYINPUT116), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n833_), .A2(new_n835_), .A3(KEYINPUT118), .A4(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n833_), .B2(new_n835_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n642_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n841_), .B2(new_n642_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n828_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT119), .B(new_n804_), .C1(new_n846_), .C2(new_n680_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n818_), .A2(new_n820_), .A3(KEYINPUT116), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n829_), .A2(KEYINPUT116), .A3(new_n819_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n834_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT117), .B(new_n643_), .C1(new_n853_), .C2(KEYINPUT58), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n854_), .A2(new_n845_), .A3(new_n839_), .A4(new_n838_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n827_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n823_), .B2(new_n640_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n680_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n802_), .A2(new_n803_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n848_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n688_), .A2(new_n490_), .A3(new_n491_), .A4(new_n433_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n847_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n423_), .A3(new_n611_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n611_), .B(KEYINPUT80), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n804_), .B1(new_n846_), .B2(new_n703_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n868_));
  AND2_X1   g667(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n867_), .B(new_n862_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n863_), .A2(new_n871_), .A3(KEYINPUT59), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n863_), .B2(KEYINPUT59), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n866_), .B(new_n870_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n865_), .B1(new_n875_), .B2(new_n423_), .ZN(G1340gat));
  OAI21_X1  g675(.A(new_n421_), .B1(new_n570_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n864_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n421_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n571_), .B(new_n870_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n421_), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n864_), .A2(new_n419_), .A3(new_n703_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n680_), .B(new_n870_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n884_), .B2(new_n419_), .ZN(G1342gat));
  NOR2_X1   g684(.A1(new_n642_), .A2(new_n417_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n870_), .B(new_n886_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n417_), .B1(new_n863_), .B2(new_n640_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(KEYINPUT122), .A3(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  AND2_X1   g692(.A1(new_n847_), .A2(new_n861_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n698_), .A2(new_n688_), .A3(new_n491_), .A4(new_n710_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n681_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n235_), .ZN(G1344gat));
  OR3_X1    g697(.A1(new_n896_), .A2(KEYINPUT124), .A3(new_n570_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n896_), .B2(new_n570_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT123), .B(G148gat), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1345gat));
  NOR2_X1   g703(.A1(new_n896_), .A2(new_n672_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n896_), .B2(new_n642_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n640_), .A2(G162gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n688_), .A2(new_n458_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n490_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n867_), .A2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G169gat), .B1(new_n913_), .B2(new_n681_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n611_), .A2(new_n307_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(new_n918_));
  OAI22_X1  g717(.A1(new_n915_), .A2(new_n916_), .B1(new_n913_), .B2(new_n918_), .ZN(G1348gat));
  NOR3_X1   g718(.A1(new_n570_), .A2(new_n308_), .A3(new_n911_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n894_), .A2(new_n698_), .A3(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n308_), .B1(new_n913_), .B2(new_n570_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT126), .Z(G1349gat));
  NOR2_X1   g723(.A1(new_n911_), .A2(new_n672_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n894_), .A2(new_n698_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n913_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n680_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n330_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n926_), .A2(new_n319_), .B1(new_n927_), .B2(new_n929_), .ZN(G1350gat));
  NAND4_X1  g729(.A1(new_n927_), .A2(new_n678_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n643_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(new_n320_), .ZN(G1351gat));
  NOR4_X1   g733(.A1(new_n698_), .A2(new_n457_), .A3(new_n401_), .A4(new_n710_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n894_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n681_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n203_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n570_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n213_), .ZN(G1353gat));
  AOI21_X1  g739(.A(new_n928_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n894_), .A2(new_n935_), .A3(new_n941_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n943_), .B2(new_n945_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n936_), .B2(new_n642_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n640_), .A2(G218gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n936_), .B2(new_n950_), .ZN(G1355gat));
endmodule


