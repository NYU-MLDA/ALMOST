//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  AOI21_X1  g000(.A(KEYINPUT98), .B1(G228gat), .B2(G233gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT21), .A3(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT21), .B1(new_n203_), .B2(new_n204_), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n206_), .C1(new_n208_), .C2(KEYINPUT97), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(KEYINPUT97), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT3), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT96), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT96), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n219_), .A2(new_n223_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G155gat), .ZN(new_n228_));
  INV_X1    g027(.A(G162gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT95), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT95), .B1(G141gat), .B2(G148gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n239_), .A3(new_n231_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n220_), .A4(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n213_), .B1(new_n234_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n202_), .B1(new_n212_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n211_), .ZN(new_n246_));
  OAI22_X1  g045(.A1(new_n246_), .A2(new_n209_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n247_));
  AND3_X1   g046(.A1(KEYINPUT98), .A2(G228gat), .A3(G233gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(new_n202_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n220_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n225_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n224_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n232_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  AND4_X1   g054(.A1(new_n220_), .A2(new_n238_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n247_), .B(new_n249_), .C1(new_n257_), .C2(new_n213_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n244_), .A2(new_n245_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT99), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n234_), .A2(new_n213_), .A3(new_n242_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G22gat), .B(G50gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT28), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT100), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n244_), .A2(new_n258_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n245_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT100), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n261_), .A2(new_n272_), .A3(new_n266_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n268_), .A2(new_n259_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n259_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT100), .B(new_n265_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n281_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G113gat), .B(G120gat), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n282_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n234_), .A2(new_n242_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n292_), .A3(KEYINPUT105), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT105), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n285_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G57gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n293_), .A2(new_n295_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n300_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n300_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT22), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(G176gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT91), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n321_), .A2(KEYINPUT91), .A3(new_n322_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT88), .B(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(G183gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT23), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n324_), .A2(new_n325_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(G169gat), .B2(G176gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G169gat), .B2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT88), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G190gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(KEYINPUT89), .A4(KEYINPUT26), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G190gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT89), .B1(new_n326_), .B2(KEYINPUT26), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n335_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT90), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT90), .B(new_n335_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n329_), .A2(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n351_), .A2(new_n353_), .B1(new_n333_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n332_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT94), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT92), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n357_), .B(KEYINPUT94), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G15gat), .B(G43gat), .Z(new_n363_));
  AND3_X1   g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n356_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n349_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n337_), .A2(new_n339_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n341_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n327_), .A2(KEYINPUT25), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G183gat), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n342_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n375_), .A3(new_n340_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT90), .B1(new_n376_), .B2(new_n335_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n355_), .B1(new_n368_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n332_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n367_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n291_), .B1(new_n366_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT93), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n366_), .A2(new_n381_), .A3(new_n291_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n387_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n382_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n315_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  INV_X1    g193(.A(new_n355_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n247_), .B1(new_n396_), .B2(new_n332_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n355_), .B(KEYINPUT102), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n322_), .A2(KEYINPUT24), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n354_), .B1(new_n404_), .B2(KEYINPUT101), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT101), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n334_), .A2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n375_), .A2(new_n403_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT103), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n323_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n321_), .A2(new_n322_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n327_), .A2(new_n336_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n411_), .A2(KEYINPUT103), .B1(new_n330_), .B2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n402_), .A2(new_n408_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n401_), .B1(new_n414_), .B2(new_n212_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n397_), .A2(new_n400_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n212_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n356_), .B2(new_n212_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n416_), .B(KEYINPUT104), .C1(new_n418_), .C2(new_n400_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT18), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n355_), .A2(KEYINPUT102), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n355_), .A2(KEYINPUT102), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n408_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n410_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n401_), .B1(new_n429_), .B2(new_n247_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n380_), .B2(new_n247_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT104), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n399_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n419_), .A2(new_n424_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n424_), .B1(new_n419_), .B2(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n394_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(new_n433_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n423_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n400_), .B1(new_n397_), .B2(new_n415_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT106), .ZN(new_n440_));
  OAI22_X1  g239(.A1(new_n439_), .A2(new_n440_), .B1(new_n431_), .B2(new_n399_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT20), .B1(new_n429_), .B2(new_n247_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n380_), .B2(new_n247_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(KEYINPUT106), .A3(new_n400_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n424_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(KEYINPUT27), .A3(new_n445_), .ZN(new_n446_));
  AND4_X1   g245(.A1(new_n280_), .A2(new_n393_), .A3(new_n436_), .A4(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n434_), .A2(new_n435_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n307_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n310_), .B1(new_n449_), .B2(new_n300_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n301_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n309_), .A2(KEYINPUT33), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n302_), .A2(new_n454_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT106), .B1(new_n443_), .B2(new_n400_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n439_), .A2(new_n440_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n418_), .A2(new_n400_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n460_), .A2(new_n462_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n437_), .A2(new_n461_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n448_), .A2(new_n456_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n436_), .A2(new_n446_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n314_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n465_), .A2(new_n279_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n389_), .A2(new_n392_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n447_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT81), .B(G15gat), .ZN(new_n472_));
  INV_X1    g271(.A(G22gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT82), .B(G1gat), .Z(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G29gat), .B(G36gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT76), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n482_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n480_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n482_), .B(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT15), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n480_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n480_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n497_), .A3(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n489_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n499_), .B(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n471_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT7), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n509_), .B(new_n510_), .C1(new_n508_), .C2(new_n507_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n507_), .A2(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(KEYINPUT66), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT67), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n518_), .A2(new_n520_), .B1(new_n507_), .B2(KEYINPUT7), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G85gat), .B(G92gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(KEYINPUT68), .B2(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n522_), .B(new_n524_), .C1(KEYINPUT68), .C2(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT9), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT10), .B(G99gat), .ZN(new_n530_));
  OAI22_X1  g329(.A1(new_n529_), .A2(new_n523_), .B1(new_n530_), .B2(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n518_), .A2(new_n520_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(G85gat), .A3(G92gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n531_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n527_), .A2(new_n490_), .A3(new_n528_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n525_), .A2(new_n526_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT77), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n490_), .A4(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n527_), .A2(new_n528_), .A3(new_n538_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n494_), .A2(new_n545_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n546_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n544_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT80), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n544_), .A2(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n544_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT36), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT78), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n557_), .A2(new_n559_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT79), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n557_), .A2(new_n572_), .A3(new_n559_), .A4(new_n568_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n564_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT37), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(KEYINPUT79), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n570_), .A2(new_n571_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT86), .ZN(new_n579_));
  INV_X1    g378(.A(G231gat), .ZN(new_n580_));
  INV_X1    g379(.A(G233gat), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(KEYINPUT11), .B2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT69), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT69), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n582_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n585_), .B(KEYINPUT69), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n588_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n582_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n590_), .A3(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n593_), .A2(new_n597_), .A3(new_n480_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n480_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n579_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n496_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(new_n597_), .A3(new_n480_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT86), .A3(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n600_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT83), .B1(new_n598_), .B2(new_n599_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT83), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n602_), .A2(new_n613_), .A3(new_n603_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT85), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n612_), .A2(new_n614_), .A3(KEYINPUT85), .A4(new_n616_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n611_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT87), .ZN(new_n622_));
  XOR2_X1   g421(.A(G176gat), .B(G204gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT73), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT74), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n624_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT71), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n595_), .A2(new_n590_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n545_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT12), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT12), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n545_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n545_), .A2(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT64), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT70), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n541_), .A2(new_n590_), .A3(new_n595_), .A4(new_n528_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT70), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n633_), .A2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n641_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n631_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n648_), .A3(new_n631_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT13), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT13), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n649_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n578_), .A2(new_n622_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n504_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n314_), .A3(new_n475_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n570_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n471_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n621_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n656_), .A2(new_n503_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n315_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n660_), .A2(new_n661_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n662_), .A2(new_n668_), .A3(new_n669_), .ZN(G1324gat));
  XNOR2_X1  g469(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n664_), .A2(new_n466_), .A3(new_n666_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G8gat), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(KEYINPUT39), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n466_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n658_), .A2(G8gat), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT107), .B1(new_n673_), .B2(G8gat), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT39), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n678_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n672_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n678_), .A2(new_n683_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n678_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n671_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n691_), .ZN(G1325gat));
  OAI21_X1  g491(.A(G15gat), .B1(new_n667_), .B2(new_n470_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT110), .Z(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n658_), .A2(G15gat), .A3(new_n470_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n667_), .B2(new_n280_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n659_), .A2(new_n473_), .A3(new_n279_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1327gat));
  INV_X1    g501(.A(G29gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n471_), .B2(new_n577_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n436_), .A2(new_n446_), .A3(new_n467_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n453_), .A2(new_n455_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n419_), .A2(new_n424_), .A3(new_n433_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n452_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n438_), .A2(new_n706_), .A3(new_n707_), .A4(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n462_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n464_), .A2(new_n314_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n279_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n470_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n447_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n578_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n704_), .A2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n652_), .A2(new_n655_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n503_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n622_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n718_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n724_), .B(new_n721_), .C1(new_n704_), .C2(new_n717_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n703_), .B1(new_n726_), .B2(new_n314_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n622_), .A2(new_n663_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n656_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n504_), .A2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(G29gat), .A3(new_n315_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n730_), .A2(G36gat), .A3(new_n679_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT111), .B1(new_n726_), .B2(new_n466_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n715_), .B2(new_n578_), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT43), .B(new_n577_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n722_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n724_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n722_), .B(KEYINPUT44), .C1(new_n737_), .C2(new_n738_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(KEYINPUT111), .A3(new_n466_), .A4(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G36gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n735_), .B1(new_n736_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT46), .B(new_n735_), .C1(new_n736_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1329gat));
  INV_X1    g547(.A(G43gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n470_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n726_), .B2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n730_), .A2(G43gat), .A3(new_n470_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n753_));
  OR3_X1    g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1330gat));
  INV_X1    g555(.A(new_n730_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G50gat), .B1(new_n757_), .B2(new_n279_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n279_), .A2(G50gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n726_), .B2(new_n759_), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n715_), .A2(new_n503_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT113), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT87), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n621_), .B(new_n763_), .ZN(new_n764_));
  AND4_X1   g563(.A1(new_n656_), .A2(new_n762_), .A3(new_n577_), .A4(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n314_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n656_), .A2(new_n503_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n664_), .A2(new_n764_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n315_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n773_), .A3(new_n466_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G64gat), .B1(new_n770_), .B2(new_n679_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT48), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1333gat));
  NOR2_X1   g576(.A1(new_n470_), .A2(G71gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT115), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n765_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G71gat), .B1(new_n770_), .B2(new_n470_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n765_), .A2(new_n785_), .A3(new_n279_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G78gat), .B1(new_n770_), .B2(new_n280_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT50), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1335gat));
  NAND4_X1  g588(.A1(new_n762_), .A2(new_n656_), .A3(new_n663_), .A4(new_n622_), .ZN(new_n790_));
  INV_X1    g589(.A(G85gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n314_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n764_), .B(new_n768_), .C1(new_n704_), .C2(new_n717_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n794_), .B2(new_n314_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT116), .ZN(G1336gat));
  AND2_X1   g596(.A1(new_n794_), .A2(new_n466_), .ZN(new_n798_));
  INV_X1    g597(.A(G92gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n466_), .A2(new_n799_), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n798_), .A2(new_n799_), .B1(new_n790_), .B2(new_n800_), .ZN(G1337gat));
  AND2_X1   g600(.A1(new_n794_), .A2(new_n750_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n470_), .A2(new_n530_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n802_), .A2(new_n505_), .B1(new_n790_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g604(.A1(new_n718_), .A2(new_n279_), .A3(new_n622_), .A4(new_n769_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(G106gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n279_), .A2(new_n506_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n790_), .B2(new_n810_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1339gat));
  NAND2_X1  g612(.A1(new_n646_), .A2(new_n648_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(new_n629_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n646_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n637_), .A2(new_n643_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT119), .A3(new_n641_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n637_), .A2(new_n642_), .A3(new_n645_), .A4(KEYINPUT55), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n638_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n640_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .A4(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n629_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n629_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n720_), .B(new_n815_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n489_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n502_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n495_), .A2(new_n497_), .A3(new_n488_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n828_), .B(new_n831_), .C1(new_n653_), .C2(new_n649_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n827_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n833_), .B2(new_n570_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n835_), .B(new_n663_), .C1(new_n827_), .C2(new_n832_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n629_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT120), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n824_), .A2(new_n840_), .A3(KEYINPUT56), .A4(new_n629_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n824_), .A2(new_n629_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n839_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n815_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n578_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n621_), .B1(new_n837_), .B2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n764_), .A2(new_n503_), .A3(new_n719_), .A4(new_n577_), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n853_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT118), .B1(new_n853_), .B2(KEYINPUT54), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(KEYINPUT54), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n852_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n466_), .A2(new_n279_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n470_), .A2(new_n315_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n720_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n764_), .B1(new_n837_), .B2(new_n851_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n857_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n861_), .B(KEYINPUT121), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n849_), .A2(new_n578_), .A3(new_n850_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n720_), .A2(new_n815_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n844_), .B2(new_n838_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n832_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n570_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n835_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n570_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n665_), .B1(new_n869_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n859_), .A4(new_n860_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n868_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n720_), .B2(KEYINPUT122), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(KEYINPUT122), .B2(new_n882_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n863_), .B1(new_n881_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n719_), .B2(KEYINPUT60), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(KEYINPUT123), .B2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n862_), .B(new_n889_), .C1(KEYINPUT123), .C2(new_n887_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n719_), .B1(new_n868_), .B2(new_n880_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n886_), .ZN(G1341gat));
  AOI21_X1  g691(.A(G127gat), .B1(new_n862_), .B2(new_n764_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT124), .B(G127gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n665_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n881_), .B2(new_n895_), .ZN(G1342gat));
  AOI21_X1  g695(.A(G134gat), .B1(new_n862_), .B2(new_n663_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n578_), .A2(G134gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT125), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n881_), .B2(new_n899_), .ZN(G1343gat));
  NOR4_X1   g699(.A1(new_n466_), .A2(new_n280_), .A3(new_n750_), .A4(new_n315_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n720_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n656_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g706(.A(new_n764_), .B(new_n901_), .C1(new_n852_), .C2(new_n857_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT126), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n903_), .A2(new_n910_), .A3(new_n764_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT127), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n909_), .A2(new_n911_), .A3(new_n914_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1346gat));
  INV_X1    g717(.A(new_n903_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G162gat), .B1(new_n919_), .B2(new_n577_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n903_), .A2(new_n229_), .A3(new_n663_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n466_), .A2(new_n393_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n279_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n720_), .B(new_n924_), .C1(new_n865_), .C2(new_n857_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G169gat), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n925_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT22), .B(G169gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n928_), .B(new_n929_), .C1(new_n931_), .C2(new_n925_), .ZN(G1348gat));
  OR2_X1    g731(.A1(new_n865_), .A2(new_n857_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n933_), .A2(new_n656_), .A3(new_n924_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n858_), .A2(new_n279_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n719_), .A2(new_n923_), .A3(new_n320_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n934_), .A2(new_n320_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n924_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n938_), .A2(new_n343_), .A3(new_n665_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n622_), .A2(new_n923_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G183gat), .B1(new_n935_), .B2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n938_), .B2(new_n577_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n663_), .A2(new_n342_), .A3(new_n403_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n938_), .B2(new_n944_), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n679_), .A2(new_n750_), .A3(new_n468_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n879_), .A2(new_n720_), .A3(new_n946_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n879_), .A2(new_n656_), .A3(new_n946_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n879_), .A2(new_n946_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n665_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT63), .B(G211gat), .Z(new_n954_));
  NAND4_X1  g753(.A1(new_n879_), .A2(new_n621_), .A3(new_n946_), .A4(new_n954_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n952_), .B2(new_n577_), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n570_), .A2(G218gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n952_), .B2(new_n958_), .ZN(G1355gat));
endmodule


