//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT84), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n206_), .B2(KEYINPUT84), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT83), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n215_));
  OR2_X1    g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT82), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT81), .B1(new_n224_), .B2(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n223_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT81), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n214_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G99gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G43gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n229_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT85), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n233_), .A2(KEYINPUT85), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(KEYINPUT85), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n235_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n232_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n243_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G197gat), .B(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(G197gat), .A2(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G211gat), .B(G218gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n255_), .A2(KEYINPUT88), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n260_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n214_), .A2(new_n264_), .A3(new_n228_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT20), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n226_), .A2(new_n223_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n268_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n211_), .A2(new_n213_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n269_), .A2(new_n207_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n264_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(KEYINPUT92), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n272_), .B2(new_n264_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n267_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n266_), .B1(new_n265_), .B2(KEYINPUT20), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n252_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT18), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  AOI21_X1  g083(.A(new_n264_), .B1(new_n214_), .B2(new_n228_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n272_), .B2(new_n264_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(new_n252_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n280_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n284_), .B1(new_n280_), .B2(new_n290_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n250_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(KEYINPUT96), .A3(new_n252_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n288_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n252_), .B1(new_n296_), .B2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT96), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n278_), .A2(new_n252_), .A3(new_n279_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n280_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT27), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305_));
  INV_X1    g104(.A(G155gat), .ZN(new_n306_));
  INV_X1    g105(.A(G162gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT86), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(G155gat), .B2(G162gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G141gat), .B(G148gat), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OR3_X1    g116(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n318_), .A2(new_n322_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n305_), .B1(new_n317_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n264_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(G228gat), .A3(G233gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT89), .ZN(new_n333_));
  INV_X1    g132(.A(G78gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n264_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(G78gat), .B1(new_n337_), .B2(KEYINPUT89), .ZN(new_n338_));
  INV_X1    g137(.A(G106gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n331_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G106gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n330_), .A3(new_n340_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n317_), .A2(new_n326_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n305_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n317_), .A2(new_n326_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT28), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT90), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n354_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n343_), .A2(new_n346_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT90), .B1(new_n363_), .B2(new_n355_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n359_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n293_), .B(new_n304_), .C1(new_n362_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT98), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n343_), .A2(new_n346_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n361_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n304_), .A4(new_n293_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n249_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(KEYINPUT94), .Z(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(KEYINPUT95), .Z(new_n383_));
  NAND3_X1  g182(.A1(new_n350_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT4), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n241_), .A2(new_n347_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n242_), .A2(KEYINPUT93), .A3(new_n350_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI211_X1 g189(.A(new_n383_), .B(new_n385_), .C1(new_n390_), .C2(KEYINPUT4), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n382_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n380_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n385_), .B1(new_n390_), .B2(KEYINPUT4), .ZN(new_n394_));
  INV_X1    g193(.A(new_n383_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n392_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n379_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NOR4_X1   g199(.A1(new_n391_), .A2(new_n400_), .A3(new_n392_), .A4(new_n380_), .ZN(new_n401_));
  AOI211_X1 g200(.A(new_n382_), .B(new_n385_), .C1(new_n390_), .C2(KEYINPUT4), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n390_), .A2(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n380_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT33), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n398_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n291_), .A2(new_n292_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT32), .B(new_n284_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n289_), .A2(new_n252_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n265_), .A2(KEYINPUT20), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT91), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n411_), .A2(new_n267_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n412_), .B2(new_n252_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n284_), .A2(KEYINPUT32), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n393_), .A2(new_n398_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n406_), .A2(new_n407_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n372_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n371_), .A2(new_n399_), .A3(new_n361_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n293_), .A2(new_n304_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n416_), .A2(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n375_), .A2(new_n399_), .B1(new_n420_), .B2(new_n249_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G230gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G57gat), .B(G64gat), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n423_), .A2(KEYINPUT11), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(KEYINPUT11), .ZN(new_n425_));
  XOR2_X1   g224(.A(G71gat), .B(G78gat), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n425_), .A2(new_n426_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT9), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G85gat), .B(G92gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n430_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT10), .B(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT64), .B(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT65), .B1(new_n434_), .B2(new_n436_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n433_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT67), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT66), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  AND2_X1   g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n442_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n447_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n443_), .A2(KEYINPUT66), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT67), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n441_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n432_), .A2(KEYINPUT8), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G99gat), .A2(G106gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT7), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n455_), .A3(new_n454_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n432_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n429_), .B(new_n458_), .C1(new_n463_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT12), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n465_), .A2(new_n466_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n462_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n470_), .A2(new_n464_), .B1(new_n472_), .B2(new_n460_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n429_), .B1(new_n473_), .B2(new_n458_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n476_));
  INV_X1    g275(.A(new_n429_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n448_), .A2(new_n449_), .A3(new_n442_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT67), .B1(new_n454_), .B2(new_n455_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n462_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n467_), .B1(new_n480_), .B2(new_n459_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n458_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n476_), .B(new_n477_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n422_), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT69), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT12), .A3(new_n468_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n483_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n422_), .ZN(new_n491_));
  OR4_X1    g290(.A1(KEYINPUT68), .A2(new_n481_), .A3(new_n482_), .A4(new_n477_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n422_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(KEYINPUT68), .A3(new_n468_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n486_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G120gat), .B(G148gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT5), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n486_), .A2(new_n491_), .A3(new_n495_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(KEYINPUT13), .A3(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT75), .B(G15gat), .ZN(new_n510_));
  INV_X1    g309(.A(G22gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT76), .B(G1gat), .Z(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(G8gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT80), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n518_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n521_), .B(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n518_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n524_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G169gat), .B(G197gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n532_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n509_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n421_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n528_), .B1(new_n473_), .B2(new_n458_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n473_), .A2(new_n458_), .A3(new_n521_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n481_), .A2(new_n482_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n528_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n551_), .A2(KEYINPUT36), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n551_), .B2(new_n552_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n544_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n548_), .B(new_n555_), .C1(new_n558_), .C2(new_n547_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT37), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT74), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n554_), .B(KEYINPUT71), .ZN(new_n564_));
  INV_X1    g363(.A(new_n548_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n547_), .B1(new_n544_), .B2(new_n557_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT72), .B(new_n564_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n559_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n563_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  AOI211_X1 g377(.A(KEYINPUT74), .B(new_n573_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n571_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n429_), .B(new_n582_), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n518_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT78), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT17), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT79), .Z(new_n593_));
  OR2_X1    g392(.A1(new_n590_), .A2(KEYINPUT17), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n591_), .A3(new_n584_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n581_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n538_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n399_), .B(KEYINPUT99), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n598_), .A2(new_n514_), .A3(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n571_), .B(KEYINPUT100), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR4_X1   g403(.A1(new_n421_), .A2(new_n596_), .A3(new_n537_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n399_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n602_), .A3(new_n607_), .ZN(G1324gat));
  NAND2_X1  g407(.A1(new_n280_), .A2(new_n290_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n294_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n303_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT27), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n413_), .B2(new_n284_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n611_), .A2(new_n250_), .B1(new_n613_), .B2(new_n302_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n598_), .A2(G8gat), .A3(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n606_), .B2(new_n614_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n615_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(G1325gat));
  INV_X1    g420(.A(new_n249_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n605_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G15gat), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n598_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n245_), .A3(new_n622_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(KEYINPUT101), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  AOI21_X1  g432(.A(new_n511_), .B1(new_n605_), .B2(new_n417_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT42), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n511_), .A3(new_n417_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  INV_X1    g436(.A(new_n596_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n537_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n577_), .A2(new_n580_), .A3(KEYINPUT102), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT102), .B1(new_n577_), .B2(new_n580_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n374_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n373_), .B1(new_n614_), .B2(new_n372_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n399_), .B(new_n622_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n420_), .A2(new_n249_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n640_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n581_), .A2(new_n640_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n421_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n639_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT44), .B1(new_n652_), .B2(KEYINPUT103), .ZN(new_n655_));
  INV_X1    g454(.A(new_n639_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n581_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n577_), .A2(new_n580_), .A3(KEYINPUT102), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n660_), .B2(new_n421_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n648_), .A2(new_n640_), .A3(new_n581_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n654_), .B1(new_n655_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(G29gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n599_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n638_), .A2(new_n571_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n421_), .A2(new_n537_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(new_n399_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n666_), .A2(new_n668_), .B1(new_n667_), .B2(new_n673_), .ZN(G1328gat));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n653_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n652_), .A2(KEYINPUT103), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n419_), .B(new_n676_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n671_), .A2(new_n681_), .A3(new_n419_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n675_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n675_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n684_), .B(new_n687_), .C1(new_n679_), .C2(G36gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n666_), .B2(new_n622_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n672_), .A2(G43gat), .A3(new_n249_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G43gat), .B1(new_n695_), .B2(new_n249_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(KEYINPUT47), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1330gat));
  OAI21_X1  g498(.A(G50gat), .B1(new_n695_), .B2(new_n372_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n372_), .A2(G50gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT106), .Z(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n672_), .B2(new_n702_), .ZN(G1331gat));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n421_), .B2(new_n536_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n536_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n648_), .A2(KEYINPUT107), .A3(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(new_n708_), .A3(new_n597_), .A4(new_n508_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n704_), .B1(new_n709_), .B2(new_n599_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n596_), .A2(new_n536_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n648_), .A2(new_n508_), .A3(new_n603_), .A4(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT109), .Z(new_n715_));
  NOR2_X1   g514(.A1(new_n399_), .A2(new_n704_), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n711_), .A2(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OR3_X1    g516(.A1(new_n709_), .A2(G64gat), .A3(new_n614_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n419_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G64gat), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT48), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT48), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1333gat));
  OR3_X1    g522(.A1(new_n709_), .A2(G71gat), .A3(new_n249_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n715_), .A2(new_n622_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G71gat), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n715_), .A2(new_n417_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G78gat), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT50), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT50), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n417_), .A2(new_n334_), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n732_), .A2(new_n733_), .B1(new_n709_), .B2(new_n734_), .ZN(G1335gat));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n706_), .A2(new_n708_), .A3(new_n508_), .A4(new_n669_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n599_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n661_), .A2(new_n662_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n509_), .A2(new_n638_), .A3(new_n536_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(new_n736_), .A3(new_n399_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n739_), .A2(new_n743_), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n742_), .B2(new_n614_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n614_), .A2(G92gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n737_), .B2(new_n746_), .ZN(G1337gat));
  NAND2_X1  g546(.A1(new_n622_), .A2(new_n435_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n737_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT112), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n740_), .A2(new_n622_), .A3(new_n741_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n751_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT111), .B1(new_n751_), .B2(G99gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n750_), .B(new_n756_), .C1(new_n753_), .C2(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1338gat));
  NAND3_X1  g557(.A1(new_n740_), .A2(new_n417_), .A3(new_n741_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G106gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n417_), .A2(new_n437_), .ZN(new_n763_));
  OAI22_X1  g562(.A1(new_n761_), .A2(new_n762_), .B1(new_n737_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n764_), .B(new_n766_), .ZN(G1339gat));
  AOI211_X1 g566(.A(new_n249_), .B(new_n599_), .C1(new_n368_), .C2(new_n374_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n535_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n529_), .A2(new_n530_), .A3(new_n525_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n526_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n490_), .B1(new_n489_), .B2(new_n422_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT69), .B(new_n493_), .C1(new_n488_), .C2(new_n483_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n502_), .B1(new_n777_), .B2(new_n495_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n503_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n504_), .A2(new_n782_), .A3(new_n774_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n536_), .A2(new_n503_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n489_), .A2(KEYINPUT55), .A3(new_n422_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n489_), .A2(new_n788_), .A3(KEYINPUT55), .A4(new_n422_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n489_), .A2(new_n422_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n500_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT56), .B(new_n500_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n785_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n571_), .B1(new_n784_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n782_), .B1(new_n504_), .B2(new_n774_), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT116), .B(new_n773_), .C1(new_n501_), .C2(new_n503_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n536_), .A2(new_n503_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n797_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n486_), .A2(new_n807_), .A3(new_n491_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n790_), .B1(KEYINPUT115), .B2(new_n786_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n789_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n500_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n805_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n804_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n571_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n801_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n810_), .A2(new_n817_), .A3(KEYINPUT56), .A4(new_n500_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n818_), .A3(new_n796_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n779_), .A2(new_n773_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT58), .B1(new_n819_), .B2(new_n820_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n577_), .A2(new_n580_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n596_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n509_), .A3(new_n713_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n825_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n536_), .B(new_n768_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(KEYINPUT119), .A3(new_n835_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n768_), .B1(new_n840_), .B2(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n840_), .B2(new_n768_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n768_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(KEYINPUT59), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n707_), .A2(new_n835_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n838_), .A2(new_n839_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n571_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n800_), .B(new_n572_), .C1(new_n804_), .C2(new_n812_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n822_), .A2(new_n823_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n821_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n638_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n826_), .A2(new_n829_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n827_), .B2(new_n826_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n825_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT60), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n509_), .B2(KEYINPUT60), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n859_), .A2(new_n768_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n509_), .B(new_n843_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n860_), .ZN(G1341gat));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n859_), .A2(new_n866_), .A3(new_n638_), .A4(new_n768_), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n596_), .B(new_n843_), .C1(new_n844_), .C2(KEYINPUT59), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n866_), .ZN(G1342gat));
  XNOR2_X1  g668(.A(KEYINPUT121), .B(G134gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n823_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n859_), .A2(new_n604_), .A3(new_n768_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n845_), .A2(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1343gat));
  NOR4_X1   g673(.A1(new_n599_), .A2(new_n372_), .A3(new_n419_), .A4(new_n622_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT122), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n536_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n508_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n638_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n878_), .B2(new_n604_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n643_), .A2(G162gat), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n877_), .B(new_n887_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n604_), .B(new_n876_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n307_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n878_), .A2(G162gat), .A3(new_n643_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(G1347gat));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n825_), .A2(new_n830_), .ZN(new_n897_));
  AND4_X1   g696(.A1(new_n372_), .A2(new_n599_), .A3(new_n419_), .A4(new_n622_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(new_n536_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  OAI21_X1  g699(.A(G169gat), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n898_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(KEYINPUT124), .A3(new_n707_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n896_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n209_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n899_), .A2(new_n900_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n902_), .B2(new_n707_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n906_), .A2(KEYINPUT62), .A3(new_n907_), .A4(G169gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n904_), .A2(new_n905_), .A3(new_n908_), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n509_), .A2(new_n210_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n859_), .A2(new_n898_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n859_), .A2(new_n913_), .A3(new_n898_), .A4(new_n910_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n210_), .B1(new_n902_), .B2(new_n509_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n912_), .A2(new_n914_), .A3(new_n915_), .ZN(G1349gat));
  NOR2_X1   g715(.A1(new_n596_), .A2(new_n223_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n897_), .A2(new_n898_), .A3(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(G183gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n859_), .A2(new_n638_), .A3(new_n898_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n902_), .B2(new_n823_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n604_), .A2(new_n226_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n902_), .B2(new_n924_), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n614_), .A2(new_n418_), .A3(new_n622_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n859_), .A2(new_n536_), .A3(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g727(.A1(new_n859_), .A2(new_n508_), .A3(new_n926_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931_));
  INV_X1    g730(.A(G211gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n638_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n859_), .A2(new_n926_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n932_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1354gat));
  NAND2_X1  g736(.A1(new_n859_), .A2(new_n926_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G218gat), .B1(new_n938_), .B2(new_n823_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n604_), .A2(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n938_), .B2(new_n941_), .ZN(G1355gat));
endmodule


