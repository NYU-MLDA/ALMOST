//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G29gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G113gat), .ZN(new_n208_));
  INV_X1    g007(.A(G120gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  INV_X1    g024(.A(G155gat), .ZN(new_n226_));
  INV_X1    g025(.A(G162gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n224_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(KEYINPUT87), .B(new_n231_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n223_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(KEYINPUT88), .B(new_n223_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n231_), .B(KEYINPUT1), .ZN(new_n240_));
  AOI211_X1 g039(.A(new_n215_), .B(new_n220_), .C1(new_n240_), .C2(new_n230_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n212_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  AOI211_X1 g042(.A(KEYINPUT89), .B(new_n241_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n211_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n241_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n210_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n248_), .B(new_n250_), .C1(KEYINPUT4), .C2(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n249_), .A3(new_n247_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n206_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n247_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n250_), .B1(new_n245_), .B2(KEYINPUT4), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n252_), .B(new_n206_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G227gat), .A2(G233gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT84), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT30), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT82), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G183gat), .A3(G190gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n266_), .A3(KEYINPUT23), .ZN(new_n267_));
  INV_X1    g066(.A(G183gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n263_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(G176gat), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n276_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT83), .B1(new_n285_), .B2(new_n279_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n274_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n264_), .A2(new_n266_), .A3(new_n272_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n263_), .A2(KEYINPUT23), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n263_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n279_), .A2(KEYINPUT24), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  MUX2_X1   g094(.A(new_n294_), .B(KEYINPUT24), .S(new_n295_), .Z(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT26), .B1(new_n269_), .B2(new_n270_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G190gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G71gat), .B(G99gat), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n287_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n287_), .B2(new_n302_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G43gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n267_), .A2(new_n273_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n278_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n285_), .A2(KEYINPUT83), .A3(new_n279_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n271_), .A2(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n293_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n303_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n287_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n307_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n262_), .B1(new_n309_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n308_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n307_), .A3(new_n316_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n261_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT31), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT31), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n318_), .A2(new_n319_), .A3(new_n325_), .A4(new_n322_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n324_), .A2(new_n210_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n210_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n243_), .A2(new_n244_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR4_X1   g132(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT29), .B1(new_n243_), .B2(new_n244_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337_));
  XOR2_X1   g136(.A(G197gat), .B(G204gat), .Z(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(KEYINPUT21), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G197gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT90), .B1(new_n340_), .B2(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n342_));
  INV_X1    g141(.A(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(G197gat), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n341_), .A2(new_n344_), .B1(new_n340_), .B2(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n339_), .B1(new_n346_), .B2(KEYINPUT21), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT21), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n337_), .B1(new_n345_), .B2(KEYINPUT91), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n336_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n246_), .B2(new_n332_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(G228gat), .A3(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n335_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G22gat), .B(G50gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G106gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n353_), .B(new_n355_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n329_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n324_), .A2(new_n326_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n211_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n324_), .A2(new_n210_), .A3(new_n326_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(new_n361_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT18), .B(G64gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G92gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n287_), .A2(new_n302_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n351_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n293_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n283_), .A2(new_n284_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT92), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n381_), .B(new_n279_), .C1(new_n383_), .C2(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n300_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT26), .B(G190gat), .Z(new_n386_));
  OAI211_X1 g185(.A(new_n310_), .B(new_n296_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n380_), .B(KEYINPUT20), .C1(new_n388_), .C2(new_n351_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n351_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n351_), .A2(new_n379_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT20), .A4(new_n391_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n378_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AND4_X1   g197(.A1(KEYINPUT20), .A2(new_n394_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n398_), .B(KEYINPUT27), .C1(new_n400_), .C2(new_n377_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n393_), .A2(new_n396_), .A3(new_n378_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n404_), .B2(new_n397_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  AND4_X1   g205(.A1(new_n258_), .A2(new_n364_), .A3(new_n373_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n256_), .A2(KEYINPUT94), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n251_), .A2(new_n409_), .A3(new_n252_), .A4(new_n206_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n251_), .A2(KEYINPUT33), .A3(new_n252_), .A4(new_n206_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n404_), .B2(new_n397_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n398_), .A2(KEYINPUT93), .A3(new_n403_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n245_), .A2(new_n418_), .A3(new_n247_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n250_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n248_), .B(new_n249_), .C1(KEYINPUT4), .C2(new_n245_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n205_), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n412_), .A2(new_n413_), .A3(new_n417_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n400_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n393_), .A2(new_n396_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n425_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n426_), .B(new_n428_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n364_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n407_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G22gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G1gat), .A2(G8gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT14), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .A4(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G29gat), .ZN(new_n443_));
  INV_X1    g242(.A(G36gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G43gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G29gat), .A2(G36gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G50gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G29gat), .B(G36gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G43gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(G50gat), .B1(new_n454_), .B2(new_n448_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n442_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n450_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(G50gat), .A3(new_n448_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n457_), .A2(new_n440_), .A3(new_n458_), .A4(new_n441_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n459_), .A3(KEYINPUT77), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT15), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n452_), .A2(new_n455_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT15), .B1(new_n457_), .B2(new_n458_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n442_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n463_), .A3(new_n459_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  INV_X1    g271(.A(G169gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G197gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT79), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n466_), .A2(new_n478_), .A3(new_n471_), .A4(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n466_), .A2(new_n471_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n475_), .B(KEYINPUT78), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G85gat), .B(G92gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(KEYINPUT9), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT9), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n491_), .A2(new_n492_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n494_), .A2(new_n495_), .A3(new_n498_), .A4(new_n496_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n500_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT65), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n500_), .A2(new_n508_), .A3(KEYINPUT65), .A4(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n452_), .A2(new_n455_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT71), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT34), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n510_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n522_), .A3(new_n515_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n517_), .A2(new_n520_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G134gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n227_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT36), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n525_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT37), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n526_), .A2(new_n532_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n540_), .B(new_n533_), .C1(new_n541_), .C2(new_n537_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G57gat), .ZN(new_n544_));
  INV_X1    g343(.A(G64gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G57gat), .A2(G64gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550_));
  INV_X1    g349(.A(G71gat), .ZN(new_n551_));
  INV_X1    g350(.A(G78gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT66), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n547_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n549_), .A2(new_n557_), .A3(new_n550_), .A4(new_n553_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  XOR2_X1   g362(.A(new_n442_), .B(KEYINPUT72), .Z(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT67), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G155gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT74), .B(G127gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n565_), .A2(KEYINPUT67), .A3(new_n566_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n567_), .A2(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n567_), .A2(KEYINPUT75), .A3(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n560_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT67), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n568_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n514_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT68), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n589_), .A2(new_n590_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n591_), .A2(new_n514_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n587_), .A2(new_n510_), .A3(KEYINPUT12), .A4(new_n588_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT69), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n561_), .A2(KEYINPUT69), .A3(KEYINPUT12), .A4(new_n510_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n601_), .A2(new_n606_), .A3(new_n597_), .A4(new_n592_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n599_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n343_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n282_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT70), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(new_n612_), .A3(new_n607_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT13), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n543_), .A2(new_n586_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT76), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n484_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n431_), .B(new_n621_), .C1(new_n620_), .C2(new_n619_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n258_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n436_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n625_));
  AND2_X1   g424(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n417_), .A2(new_n423_), .A3(new_n413_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n429_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n364_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n364_), .A2(new_n373_), .A3(new_n406_), .A4(new_n258_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n585_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n534_), .A2(new_n538_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT13), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n617_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n484_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n635_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n258_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT97), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n627_), .B(new_n642_), .C1(new_n625_), .C2(new_n624_), .ZN(G1324gat));
  OAI21_X1  g442(.A(G8gat), .B1(new_n640_), .B2(new_n406_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT99), .B(KEYINPUT39), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n406_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n437_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g449(.A(G15gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n622_), .A2(new_n651_), .A3(new_n368_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G15gat), .B1(new_n640_), .B2(new_n329_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT100), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT100), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(KEYINPUT41), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n654_), .B2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n656_), .B2(new_n657_), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n362_), .A2(new_n363_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n640_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n622_), .A2(new_n663_), .A3(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1327gat));
  NOR3_X1   g464(.A1(new_n637_), .A2(new_n586_), .A3(new_n638_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n539_), .A2(new_n542_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n407_), .B2(new_n430_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n632_), .A2(new_n633_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n668_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n667_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n674_), .B2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n671_), .B2(new_n668_), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT43), .B(new_n543_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n666_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(KEYINPUT44), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n623_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n635_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n666_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n258_), .A2(G29gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT102), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n684_), .A2(new_n443_), .B1(new_n687_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT104), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT104), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n406_), .B1(new_n674_), .B2(KEYINPUT44), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n444_), .B1(new_n682_), .B2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n685_), .A2(new_n444_), .A3(new_n666_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n696_), .A2(KEYINPUT103), .A3(new_n406_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT103), .B1(new_n696_), .B2(new_n406_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n692_), .B(new_n693_), .C1(new_n695_), .C2(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n674_), .A2(KEYINPUT101), .A3(KEYINPUT44), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n694_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n698_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n698_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n708_), .A2(KEYINPUT104), .A3(new_n691_), .A4(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n704_), .A2(new_n712_), .ZN(G1329gat));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n368_), .B(new_n683_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G43gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n329_), .A2(G43gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n686_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT47), .B(new_n720_), .C1(new_n715_), .C2(G43gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  NAND4_X1  g521(.A1(new_n682_), .A2(G50gat), .A3(new_n659_), .A4(new_n683_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G50gat), .B1(new_n686_), .B2(new_n659_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT105), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n728_), .A3(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n618_), .A2(new_n484_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n634_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n635_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G57gat), .A3(new_n623_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n732_), .A2(new_n668_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n623_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n544_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT106), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT106), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT107), .ZN(G1332gat));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n545_), .A3(new_n647_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n734_), .A2(new_n647_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G64gat), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT48), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(KEYINPUT48), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT108), .ZN(G1333gat));
  AOI21_X1  g548(.A(new_n551_), .B1(new_n734_), .B2(new_n368_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n551_), .A3(new_n368_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n659_), .A2(new_n552_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT110), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n736_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n552_), .B1(new_n734_), .B2(new_n659_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n758_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(KEYINPUT50), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n759_), .B2(new_n760_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n731_), .A2(new_n585_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n431_), .A2(new_n764_), .A3(new_n635_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n623_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT111), .Z(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n258_), .A2(new_n504_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(G1336gat));
  AOI21_X1  g569(.A(G92gat), .B1(new_n765_), .B2(new_n647_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n406_), .A2(new_n505_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n768_), .B2(new_n772_), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n501_), .A3(new_n368_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n768_), .A2(new_n368_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G99gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT112), .B(new_n486_), .C1(new_n768_), .C2(new_n368_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT113), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n779_), .B(new_n781_), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n765_), .A2(new_n487_), .A3(new_n659_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n659_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(G106gat), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT52), .B(new_n487_), .C1(new_n768_), .C2(new_n659_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g588(.A1(new_n616_), .A2(new_n484_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT115), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n616_), .A2(new_n484_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n601_), .A2(new_n592_), .A3(new_n606_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n598_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n607_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n796_), .A2(new_n795_), .A3(new_n598_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n614_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n589_), .A2(new_n590_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n600_), .B2(new_n594_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n597_), .B1(new_n805_), .B2(new_n606_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n607_), .B1(new_n806_), .B2(new_n795_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n800_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n794_), .B1(new_n803_), .B2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n812_), .A2(KEYINPUT116), .A3(new_n475_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n470_), .A2(new_n464_), .A3(new_n459_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT116), .B1(new_n812_), .B2(new_n475_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n813_), .A2(KEYINPUT117), .A3(new_n814_), .A4(new_n815_), .ZN(new_n819_));
  AND4_X1   g618(.A1(new_n617_), .A2(new_n480_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n635_), .B1(new_n811_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT57), .B(new_n635_), .C1(new_n811_), .C2(new_n820_), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n616_), .A2(new_n818_), .A3(new_n480_), .A4(new_n819_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n614_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n802_), .B(new_n613_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n825_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n668_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n823_), .A2(new_n824_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n585_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n619_), .B2(new_n484_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n637_), .A2(new_n668_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(new_n586_), .A3(new_n638_), .A4(new_n835_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n659_), .B1(new_n834_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n647_), .A2(new_n258_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n368_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n484_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n841_), .A2(KEYINPUT59), .A3(new_n368_), .A4(new_n842_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n638_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g649(.A(new_n209_), .B1(new_n618_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n844_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n209_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n618_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n209_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n844_), .B2(new_n586_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n848_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n586_), .A2(G127gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT118), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n856_), .B2(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n844_), .B2(new_n733_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n668_), .A2(G134gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT119), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n856_), .B2(new_n862_), .ZN(G1343gat));
  AOI211_X1 g662(.A(new_n368_), .B(new_n660_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n842_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n834_), .A2(new_n840_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n329_), .A3(new_n659_), .A4(new_n842_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n484_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G141gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n864_), .A2(KEYINPUT120), .A3(new_n842_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n213_), .A3(new_n484_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(G1344gat));
  XNOR2_X1  g675(.A(KEYINPUT121), .B(G148gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(new_n637_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n877_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n618_), .B(new_n879_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n874_), .B2(new_n586_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n882_), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n585_), .B(new_n884_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n874_), .B2(new_n733_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n227_), .B(new_n543_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n623_), .A2(new_n406_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n638_), .A2(new_n383_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n841_), .A2(new_n368_), .A3(new_n890_), .A4(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n484_), .A3(new_n368_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT122), .ZN(new_n894_));
  AOI211_X1 g693(.A(KEYINPUT62), .B(new_n473_), .C1(new_n841_), .C2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n866_), .A2(new_n660_), .A3(new_n894_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(G169gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n892_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT123), .B(new_n892_), .C1(new_n895_), .C2(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1348gat));
  NAND3_X1  g702(.A1(new_n841_), .A2(new_n368_), .A3(new_n890_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n618_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n282_), .ZN(G1349gat));
  OAI21_X1  g705(.A(G183gat), .B1(new_n904_), .B2(new_n585_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n904_), .A2(new_n585_), .A3(new_n385_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT124), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  OR3_X1    g709(.A1(new_n904_), .A2(new_n585_), .A3(new_n385_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n907_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n904_), .B2(new_n543_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n635_), .A2(new_n386_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n904_), .B2(new_n916_), .ZN(G1351gat));
  AND2_X1   g716(.A1(new_n864_), .A2(new_n890_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n918_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n484_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n864_), .A2(new_n484_), .A3(new_n890_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n340_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n920_), .B2(new_n340_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n919_), .A2(new_n921_), .A3(new_n923_), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n864_), .A2(new_n890_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n618_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n343_), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n864_), .A2(new_n586_), .A3(new_n890_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(KEYINPUT127), .A3(new_n929_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT63), .B(G211gat), .Z(new_n934_));
  NAND4_X1  g733(.A1(new_n918_), .A2(KEYINPUT126), .A3(new_n586_), .A4(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  INV_X1    g735(.A(new_n934_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n928_), .B2(new_n937_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n932_), .A2(new_n933_), .B1(new_n935_), .B2(new_n938_), .ZN(G1354gat));
  AOI21_X1  g738(.A(G218gat), .B1(new_n918_), .B2(new_n733_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n925_), .A2(new_n543_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(G218gat), .B2(new_n941_), .ZN(G1355gat));
endmodule


