//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT87), .B(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n211_), .A2(KEYINPUT88), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT88), .B2(new_n211_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT24), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n213_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n230_), .A2(KEYINPUT92), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT92), .B1(new_n230_), .B2(new_n231_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n231_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n233_), .A2(KEYINPUT93), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(KEYINPUT93), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n230_), .A2(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n206_), .B1(new_n229_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT25), .B(G183gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n219_), .A2(new_n243_), .B1(new_n244_), .B2(new_n224_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n225_), .A2(new_n210_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n245_), .B(new_n213_), .C1(new_n246_), .C2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n210_), .A2(KEYINPUT98), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n210_), .A2(KEYINPUT98), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n248_), .A2(new_n209_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n251_), .A3(new_n236_), .A4(new_n240_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT99), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n242_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G8gat), .B(G36gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n218_), .A2(new_n240_), .A3(new_n236_), .A4(new_n228_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(new_n247_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n204_), .B1(new_n263_), .B2(new_n241_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n203_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT27), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n261_), .B(KEYINPUT104), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n203_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n203_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n252_), .A2(KEYINPUT20), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n229_), .A2(new_n241_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n269_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT105), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT105), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(new_n269_), .C1(new_n270_), .C2(new_n274_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n268_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT102), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n252_), .B(new_n253_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n281_), .A2(new_n242_), .B1(new_n265_), .B2(new_n203_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n282_), .B2(new_n261_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n256_), .A2(new_n266_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n261_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT102), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT101), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n282_), .B2(new_n261_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AND4_X1   g089(.A1(new_n288_), .A2(new_n256_), .A3(new_n261_), .A4(new_n266_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n279_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(G127gat), .B(G134gat), .Z(new_n297_));
  XOR2_X1   g096(.A(G113gat), .B(G120gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OR3_X1    g099(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT90), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n312_), .A3(new_n309_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G141gat), .ZN(new_n315_));
  INV_X1    g114(.A(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n308_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n302_), .B(new_n317_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n300_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n299_), .A2(new_n314_), .A3(new_n321_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT4), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n300_), .A2(new_n326_), .A3(new_n322_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n296_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n296_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n328_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n333_), .B1(new_n328_), .B2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n241_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n342_), .A2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n340_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n340_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n345_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT94), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT95), .B(new_n340_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n351_), .A2(new_n356_), .A3(new_n345_), .A4(new_n352_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n350_), .A2(new_n354_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n353_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n353_), .A2(new_n366_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n363_), .A3(new_n348_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT31), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n229_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n299_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n299_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n377_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n295_), .A2(new_n339_), .A3(new_n371_), .A4(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n338_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n289_), .A2(new_n291_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n325_), .A2(new_n296_), .A3(new_n327_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n323_), .A2(new_n334_), .A3(new_n324_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT103), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n332_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n393_), .B2(new_n332_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n337_), .A2(KEYINPUT33), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n333_), .C1(new_n328_), .C2(new_n335_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n402_), .A3(new_n287_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n261_), .A2(KEYINPUT32), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n338_), .B(new_n405_), .C1(new_n284_), .C2(new_n404_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n390_), .A2(new_n295_), .B1(new_n407_), .B2(new_n371_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n387_), .B(KEYINPUT89), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n389_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT107), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT66), .B(G85gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT9), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(G92gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n415_));
  OR2_X1    g214(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT9), .A3(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n414_), .A2(new_n419_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT67), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n422_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT67), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n419_), .A4(new_n414_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G29gat), .B(G36gat), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT74), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(KEYINPUT74), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G43gat), .B(G50gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT68), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n447_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n420_), .A2(KEYINPUT69), .A3(new_n421_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n456_));
  AND2_X1   g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT8), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n441_), .B1(new_n454_), .B2(new_n461_), .ZN(new_n462_));
  NOR4_X1   g261(.A1(KEYINPUT68), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n452_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n425_), .B(new_n446_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n455_), .A2(new_n459_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT70), .A4(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n443_), .A2(KEYINPUT71), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT71), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT6), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n442_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n446_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n451_), .A2(new_n453_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n471_), .A3(new_n442_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n460_), .B1(new_n477_), .B2(new_n466_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n431_), .B(new_n440_), .C1(new_n468_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT75), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n455_), .A2(new_n459_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n469_), .A2(new_n471_), .A3(new_n442_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n482_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(new_n475_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n462_), .B(new_n467_), .C1(new_n484_), .C2(new_n460_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT75), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n431_), .A4(new_n440_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT78), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n490_));
  AND2_X1   g289(.A1(G232gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT35), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n438_), .A2(KEYINPUT15), .A3(new_n439_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT15), .B1(new_n438_), .B2(new_n439_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n431_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n488_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n489_), .B1(new_n488_), .B2(new_n498_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(KEYINPUT35), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n480_), .A2(new_n487_), .B1(new_n497_), .B2(new_n496_), .ZN(new_n502_));
  OAI22_X1  g301(.A1(new_n499_), .A2(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G190gat), .B(G218gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT76), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n499_), .A2(new_n500_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT77), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n496_), .A2(new_n497_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n488_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n501_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n503_), .A2(KEYINPUT80), .A3(new_n508_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n410_), .A2(new_n411_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n411_), .B1(new_n410_), .B2(new_n523_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G57gat), .B(G64gat), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n530_));
  XOR2_X1   g329(.A(G71gat), .B(G78gat), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n431_), .B(new_n534_), .C1(new_n468_), .C2(new_n478_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT64), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  INV_X1    g339(.A(new_n534_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n497_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n497_), .B2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n534_), .B1(new_n485_), .B2(new_n431_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n535_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n537_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT72), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT81), .B(G1gat), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n561_), .A2(G8gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT14), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G1gat), .B(G8gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n496_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n440_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n566_), .A2(new_n568_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT86), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT85), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n572_), .A2(new_n575_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n555_), .A2(KEYINPUT13), .A3(new_n556_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n559_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT106), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n559_), .A2(KEYINPUT106), .A3(new_n584_), .A4(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n534_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n566_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT84), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT82), .A3(KEYINPUT17), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n594_), .B(new_n601_), .C1(KEYINPUT17), .C2(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n591_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n527_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n338_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G1gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT27), .B1(new_n391_), .B2(new_n287_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n386_), .A2(new_n384_), .A3(new_n339_), .ZN(new_n610_));
  NOR4_X1   g409(.A1(new_n609_), .A2(new_n370_), .A3(new_n610_), .A4(new_n279_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n407_), .A2(new_n371_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n293_), .A2(new_n294_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n279_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n390_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n409_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n586_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n503_), .A2(KEYINPUT80), .A3(new_n508_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT80), .B1(new_n503_), .B2(new_n508_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT37), .B1(new_n512_), .B2(new_n520_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT79), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n499_), .A2(new_n500_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n516_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n502_), .B2(new_n501_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n520_), .B(KEYINPUT79), .C1(new_n500_), .C2(new_n499_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n509_), .A3(new_n629_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n622_), .A2(new_n623_), .B1(new_n630_), .B2(KEYINPUT37), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n604_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n619_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n339_), .A2(new_n561_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n608_), .A2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(G8gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n295_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n639_), .B(new_n605_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  AND4_X1   g441(.A1(KEYINPUT108), .A2(new_n641_), .A3(new_n642_), .A4(G8gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT108), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n638_), .B1(new_n644_), .B2(KEYINPUT39), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n641_), .A2(new_n645_), .B1(KEYINPUT108), .B2(new_n642_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n640_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1325gat));
  NAND3_X1  g448(.A1(new_n633_), .A2(new_n373_), .A3(new_n409_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n606_), .A2(new_n409_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT41), .B1(new_n651_), .B2(G15gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n633_), .A2(new_n655_), .A3(new_n370_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n606_), .A2(new_n370_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G22gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT42), .B(new_n655_), .C1(new_n606_), .C2(new_n370_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1327gat));
  XOR2_X1   g460(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n662_));
  NAND2_X1  g461(.A1(new_n630_), .A2(KEYINPUT37), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n511_), .A2(new_n522_), .A3(new_n623_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n618_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n410_), .A2(new_n631_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n590_), .A2(new_n604_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n672_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(new_n338_), .ZN(new_n678_));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n604_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n523_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n619_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n338_), .A2(new_n679_), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n678_), .A2(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  OR3_X1    g483(.A1(new_n682_), .A2(G36gat), .A3(new_n295_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT45), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n676_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT44), .B(new_n672_), .C1(new_n666_), .C2(new_n669_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n687_), .B(new_n639_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n677_), .B2(new_n639_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n686_), .B(KEYINPUT46), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n677_), .B2(new_n388_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n682_), .A2(G43gat), .A3(new_n617_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n701_));
  OR3_X1    g500(.A1(new_n699_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1330gat));
  OR3_X1    g503(.A1(new_n682_), .A2(G50gat), .A3(new_n371_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n677_), .A2(new_n370_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT113), .B1(new_n706_), .B2(G50gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1331gat));
  AND2_X1   g508(.A1(new_n559_), .A2(new_n585_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n584_), .A2(new_n604_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n527_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(G57gat), .A3(new_n338_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT115), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT115), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n631_), .A2(new_n710_), .A3(new_n604_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(KEYINPUT114), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n618_), .A2(new_n584_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(KEYINPUT114), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n338_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n715_), .A2(new_n716_), .A3(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n725_), .A3(new_n639_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n713_), .A2(new_n639_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G64gat), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT48), .B(new_n725_), .C1(new_n713_), .C2(new_n639_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n732_), .A3(new_n409_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n713_), .A2(new_n409_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G71gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT49), .B(new_n732_), .C1(new_n713_), .C2(new_n409_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n722_), .A2(new_n739_), .A3(new_n370_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n713_), .A2(new_n370_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n739_), .C1(new_n713_), .C2(new_n370_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  AND3_X1   g544(.A1(new_n719_), .A2(new_n711_), .A3(new_n681_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n338_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n582_), .A2(new_n583_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n711_), .A2(new_n604_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n338_), .A2(new_n412_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT116), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n750_), .B2(new_n752_), .ZN(G1336gat));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n754_), .A3(new_n639_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n750_), .A2(new_n639_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n754_), .ZN(G1337gat));
  NAND4_X1  g556(.A1(new_n746_), .A2(new_n415_), .A3(new_n417_), .A4(new_n388_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n409_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G99gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G99gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(KEYINPUT118), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n763_), .B(new_n765_), .ZN(G1338gat));
  NAND4_X1  g565(.A1(new_n746_), .A2(new_n416_), .A3(new_n418_), .A4(new_n370_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n370_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g572(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n710_), .A2(new_n665_), .A3(new_n712_), .A4(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n710_), .A2(new_n665_), .A3(new_n712_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n535_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n537_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n544_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT55), .B(new_n539_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n552_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n548_), .A2(new_n553_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n567_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n571_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n579_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n572_), .A2(new_n575_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n580_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n792_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n780_), .B1(new_n791_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT121), .B1(new_n801_), .B2(new_n665_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n552_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n779_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n631_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n800_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n802_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n584_), .A2(new_n792_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n555_), .A2(new_n556_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT57), .B(new_n523_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n748_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n557_), .A2(new_n799_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n819_), .B2(new_n523_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n810_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n778_), .B1(new_n822_), .B2(new_n604_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n639_), .A2(new_n370_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n338_), .A3(new_n388_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n825_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n680_), .B1(new_n810_), .B2(new_n821_), .ZN(new_n832_));
  OAI221_X1 g631(.A(new_n830_), .B1(new_n831_), .B2(new_n828_), .C1(new_n832_), .C2(new_n778_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n584_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G113gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n826_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n748_), .A2(G113gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(G1340gat));
  AND3_X1   g637(.A1(new_n829_), .A2(new_n711_), .A3(new_n833_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n710_), .B2(KEYINPUT60), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(KEYINPUT60), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(KEYINPUT123), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(KEYINPUT123), .B2(new_n841_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n839_), .A2(new_n840_), .B1(new_n836_), .B2(new_n844_), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n829_), .A2(new_n680_), .A3(new_n833_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G127gat), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n604_), .A2(G127gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n836_), .B2(new_n848_), .ZN(G1342gat));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n836_), .B2(new_n523_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n665_), .A2(new_n850_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n833_), .B(new_n852_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n851_), .A2(KEYINPUT124), .A3(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1343gat));
  NAND3_X1  g657(.A1(new_n617_), .A2(new_n338_), .A3(new_n370_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n823_), .A2(new_n639_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n584_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n711_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n680_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n523_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n860_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n860_), .A2(new_n631_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(new_n868_), .ZN(G1347gat));
  NOR3_X1   g672(.A1(new_n617_), .A2(new_n338_), .A3(new_n295_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n371_), .B(new_n874_), .C1(new_n832_), .C2(new_n778_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875_), .B2(new_n748_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT125), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(G169gat), .C1(new_n875_), .C2(new_n748_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(KEYINPUT62), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n207_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n823_), .A2(new_n370_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n584_), .A3(new_n874_), .ZN(new_n883_));
  OAI221_X1 g682(.A(new_n880_), .B1(KEYINPUT62), .B2(new_n877_), .C1(new_n881_), .C2(new_n883_), .ZN(G1348gat));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n823_), .B2(new_n370_), .ZN(new_n886_));
  OAI211_X1 g685(.A(KEYINPUT126), .B(new_n371_), .C1(new_n832_), .C2(new_n778_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n874_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(new_n208_), .A3(new_n710_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n882_), .A2(new_n711_), .A3(new_n874_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n888_), .A2(new_n890_), .B1(new_n208_), .B2(new_n891_), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n604_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n887_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n214_), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n875_), .A2(new_n243_), .A3(new_n604_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT127), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n896_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n875_), .B2(new_n665_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n869_), .A2(new_n219_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n875_), .B2(new_n903_), .ZN(G1351gat));
  INV_X1    g703(.A(new_n823_), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n409_), .A2(new_n295_), .A3(new_n338_), .A4(new_n371_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n584_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n711_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  NOR4_X1   g713(.A1(new_n907_), .A2(new_n604_), .A3(new_n913_), .A4(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n908_), .A2(new_n680_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n913_), .ZN(G1354gat));
  OAI21_X1  g716(.A(G218gat), .B1(new_n907_), .B2(new_n665_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n523_), .A2(G218gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n907_), .B2(new_n919_), .ZN(G1355gat));
endmodule


