//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT97), .B1(new_n205_), .B2(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT100), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(KEYINPUT21), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT101), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT101), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT24), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n227_), .A2(new_n231_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n232_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(KEYINPUT89), .A2(G169gat), .A3(G176gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n224_), .B(new_n226_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n222_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n217_), .A2(new_n239_), .A3(new_n218_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT102), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n217_), .A2(new_n239_), .A3(KEYINPUT102), .A4(new_n218_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G169gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT99), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n210_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n208_), .A2(new_n204_), .A3(new_n250_), .A4(new_n206_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(KEYINPUT98), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT98), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n207_), .A2(new_n254_), .A3(new_n250_), .A4(new_n208_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(KEYINPUT98), .ZN(new_n257_));
  INV_X1    g056(.A(new_n251_), .ZN(new_n258_));
  AND4_X1   g057(.A1(new_n248_), .A2(new_n255_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n214_), .B(new_n247_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT103), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT103), .ZN(new_n262_));
  INV_X1    g061(.A(new_n214_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n258_), .A3(new_n257_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT99), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n248_), .A3(new_n255_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n267_), .B2(new_n247_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n223_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n219_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT24), .B1(new_n231_), .B2(new_n232_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT90), .B1(new_n277_), .B2(new_n219_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n232_), .A4(new_n233_), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT88), .B1(new_n280_), .B2(KEYINPUT25), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n221_), .B(new_n281_), .C1(new_n220_), .C2(KEYINPUT88), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .A4(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n245_), .A2(new_n240_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT20), .B(new_n272_), .C1(new_n288_), .C2(new_n267_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT104), .B1(new_n269_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n260_), .A2(KEYINPUT103), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n267_), .A2(new_n262_), .A3(new_n247_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n283_), .A2(new_n285_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n214_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n294_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT104), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n293_), .A2(new_n300_), .A3(new_n301_), .A4(new_n272_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n290_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n294_), .B1(new_n288_), .B2(new_n267_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n267_), .A2(new_n247_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n272_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G8gat), .B(G36gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT18), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n303_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n304_), .A2(new_n272_), .A3(new_n305_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n272_), .B1(new_n300_), .B2(new_n260_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(KEYINPUT27), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n311_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n320_));
  AOI211_X1 g119(.A(new_n313_), .B(new_n306_), .C1(new_n290_), .C2(new_n302_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT107), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT107), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n324_), .B(new_n319_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n318_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT0), .B(G57gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  OR2_X1    g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT95), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n343_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT2), .Z(new_n348_));
  OAI211_X1 g147(.A(new_n339_), .B(new_n340_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n340_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n343_), .B(new_n347_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n338_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n336_), .A2(new_n337_), .A3(new_n349_), .A4(new_n353_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT4), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n338_), .A2(new_n358_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n331_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n367_), .A2(new_n330_), .A3(new_n364_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G71gat), .B(G99gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT92), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT30), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n298_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(G15gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n378_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT31), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT31), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n338_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n383_), .A2(new_n337_), .A3(new_n336_), .A4(new_n385_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n370_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G22gat), .B(G50gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(new_n354_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n299_), .B(new_n394_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n394_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n395_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n267_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT28), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n402_), .A2(new_n404_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n391_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n391_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n326_), .A2(new_n389_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT32), .B(new_n311_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT106), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n369_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n413_), .A2(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n311_), .A2(KEYINPUT32), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n303_), .A2(new_n307_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n303_), .A2(new_n307_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n313_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT105), .B1(new_n366_), .B2(KEYINPUT33), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n330_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT105), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n357_), .A2(new_n361_), .A3(new_n359_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n355_), .A2(new_n356_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n330_), .B1(new_n430_), .B2(new_n362_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n366_), .A2(KEYINPUT33), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n421_), .A2(new_n427_), .A3(new_n312_), .A4(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n412_), .B1(new_n419_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n369_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n326_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n387_), .A2(new_n388_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n411_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT6), .Z(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  INV_X1    g241(.A(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G106gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT67), .B1(new_n441_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n440_), .B(KEYINPUT6), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n446_), .A4(new_n445_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G85gat), .B(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n447_), .B1(new_n449_), .B2(new_n455_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G92gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(KEYINPUT9), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n461_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT9), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n441_), .B1(new_n468_), .B2(KEYINPUT66), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT64), .B(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(KEYINPUT65), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n460_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n483_));
  XOR2_X1   g282(.A(G71gat), .B(G78gat), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT12), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT72), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n472_), .A2(KEYINPUT65), .A3(new_n473_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT65), .B1(new_n472_), .B2(new_n473_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n471_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n467_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n464_), .A2(new_n466_), .B1(new_n465_), .B2(G92gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT66), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n449_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n491_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n469_), .A2(KEYINPUT71), .A3(new_n478_), .A4(new_n471_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n460_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n488_), .ZN(new_n502_));
  AND2_X1   g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n460_), .A2(new_n479_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(new_n487_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n490_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT73), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n487_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT70), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n480_), .A2(new_n488_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n503_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n490_), .A2(new_n513_), .A3(new_n502_), .A4(new_n505_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G120gat), .B(G148gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G176gat), .B(G204gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n507_), .A2(new_n512_), .A3(new_n514_), .A4(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT78), .B(G1gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT79), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G8gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n532_), .B(KEYINPUT79), .ZN(new_n537_));
  INV_X1    g336(.A(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G29gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n536_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(G229gat), .A3(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n543_), .B(KEYINPUT15), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT84), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT84), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n546_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT85), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n548_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT87), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT86), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n557_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n527_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n439_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G127gat), .B(G155gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n540_), .B(KEYINPUT81), .ZN(new_n574_));
  AND2_X1   g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n487_), .B(KEYINPUT80), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n573_), .B1(new_n578_), .B2(KEYINPUT83), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n573_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(KEYINPUT17), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n579_), .A2(KEYINPUT17), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT77), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n504_), .A2(new_n543_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n501_), .A2(KEYINPUT75), .A3(new_n549_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT75), .B1(new_n501_), .B2(new_n549_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT76), .B1(new_n597_), .B2(new_n598_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n594_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n594_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n589_), .B(new_n591_), .C1(new_n603_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n598_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n501_), .A2(KEYINPUT75), .A3(new_n549_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n600_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n602_), .A3(new_n595_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT35), .A3(new_n593_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n606_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n588_), .A3(new_n587_), .A4(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n614_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n583_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n567_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n370_), .A3(new_n528_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT38), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n607_), .A2(new_n614_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n583_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n567_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(new_n369_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(new_n326_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n621_), .A2(new_n529_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(new_n627_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n630_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n634_), .B2(G8gat), .ZN(new_n635_));
  AOI211_X1 g434(.A(KEYINPUT39), .B(new_n529_), .C1(new_n633_), .C2(new_n630_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(new_n438_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n627_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n621_), .A2(new_n377_), .A3(new_n438_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  OAI21_X1  g444(.A(G22gat), .B1(new_n627_), .B2(new_n410_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT42), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n410_), .A2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n620_), .B2(new_n648_), .ZN(G1327gat));
  OR2_X1    g448(.A1(new_n581_), .A2(new_n582_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n624_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n567_), .A2(new_n651_), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n652_), .A2(G29gat), .A3(new_n369_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n439_), .A2(new_n655_), .A3(new_n618_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT37), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n624_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n614_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(KEYINPUT109), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n435_), .B(new_n318_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n640_), .B1(new_n665_), .B2(new_n434_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(new_n411_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT110), .B1(new_n667_), .B2(new_n655_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n659_), .A2(new_n663_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n421_), .A2(new_n312_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n324_), .B1(new_n670_), .B2(new_n319_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n325_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n436_), .B(new_n317_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n434_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n438_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n326_), .A2(new_n389_), .A3(new_n410_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(KEYINPUT43), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n657_), .B1(new_n668_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n566_), .A2(new_n583_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n654_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT110), .B(new_n655_), .C1(new_n439_), .C2(new_n669_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n677_), .B2(KEYINPUT43), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n656_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n681_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n370_), .A3(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT111), .A3(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT111), .B1(new_n688_), .B2(G29gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n653_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n630_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n652_), .A2(G36gat), .A3(new_n326_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT45), .Z(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n695_), .A3(KEYINPUT46), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n682_), .A2(new_n687_), .A3(G43gat), .A4(new_n438_), .ZN(new_n701_));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n652_), .B2(new_n640_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1330gat));
  AND2_X1   g505(.A1(new_n682_), .A2(new_n687_), .ZN(new_n707_));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n410_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n567_), .A2(new_n412_), .A3(new_n651_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n707_), .A2(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(G1331gat));
  AND3_X1   g510(.A1(new_n439_), .A2(new_n565_), .A3(new_n527_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n626_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n369_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n619_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n369_), .A2(G57gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n713_), .B2(new_n326_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n326_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n715_), .B2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n713_), .B2(new_n640_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n640_), .A2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n715_), .B2(new_n724_), .ZN(G1334gat));
  OR3_X1    g524(.A1(new_n715_), .A2(G78gat), .A3(new_n410_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G78gat), .B1(new_n713_), .B2(new_n410_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT113), .Z(G1335gat));
  NAND2_X1  g530(.A1(new_n712_), .A2(new_n651_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n463_), .A3(new_n370_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n527_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n650_), .A2(new_n736_), .A3(new_n564_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n685_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n370_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n739_), .B2(new_n463_), .ZN(G1336gat));
  NOR2_X1   g539(.A1(new_n326_), .A2(new_n461_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT115), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G92gat), .B1(new_n734_), .B2(new_n630_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1337gat));
  AND2_X1   g547(.A1(new_n438_), .A2(new_n472_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n734_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n443_), .B1(new_n738_), .B2(new_n438_), .ZN(new_n751_));
  OR3_X1    g550(.A1(new_n750_), .A2(new_n751_), .A3(KEYINPUT51), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT51), .B1(new_n750_), .B2(new_n751_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n734_), .A2(new_n473_), .A3(new_n412_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n685_), .A2(new_n412_), .A3(new_n737_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n755_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  NOR3_X1   g563(.A1(new_n630_), .A2(new_n369_), .A3(new_n412_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n547_), .A2(new_n556_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n767_));
  MUX2_X1   g566(.A(new_n767_), .B(new_n557_), .S(new_n561_), .Z(new_n768_));
  NAND2_X1  g567(.A1(new_n524_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT118), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n524_), .A2(new_n771_), .A3(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n564_), .A2(new_n523_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n507_), .A2(new_n775_), .A3(new_n514_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n509_), .A2(new_n490_), .A3(new_n502_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n503_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n775_), .B2(new_n506_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n521_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT56), .B(new_n521_), .C1(new_n777_), .C2(new_n780_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n774_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n624_), .B1(new_n773_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI221_X1 g587(.A(new_n624_), .B1(KEYINPUT119), .B2(KEYINPUT57), .C1(new_n773_), .C2(new_n785_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n776_), .B(new_n779_), .C1(new_n775_), .C2(new_n506_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n521_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n794_), .A3(new_n783_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n768_), .A2(new_n523_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(KEYINPUT58), .A3(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n618_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n650_), .B1(new_n790_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n650_), .A2(new_n617_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n736_), .A2(new_n565_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n803_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n619_), .A2(new_n565_), .A3(new_n736_), .A4(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n438_), .B(new_n765_), .C1(new_n802_), .C2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n789_), .A3(new_n788_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n583_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n815_), .A2(new_n438_), .A3(new_n765_), .A4(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n812_), .A2(new_n818_), .A3(new_n564_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G113gat), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n810_), .A2(G113gat), .A3(new_n565_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1340gat));
  NAND3_X1  g621(.A1(new_n812_), .A2(new_n818_), .A3(new_n527_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G120gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n809_), .B1(new_n813_), .B2(new_n583_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n640_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n736_), .A2(KEYINPUT60), .ZN(new_n827_));
  MUX2_X1   g626(.A(new_n827_), .B(KEYINPUT60), .S(G120gat), .Z(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n765_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(G1341gat));
  OR2_X1    g629(.A1(KEYINPUT122), .A2(G127gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(G127gat), .B1(new_n583_), .B2(KEYINPUT122), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n812_), .A2(new_n818_), .A3(new_n831_), .A4(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n810_), .B2(new_n583_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1342gat));
  NAND3_X1  g635(.A1(new_n812_), .A2(new_n818_), .A3(new_n618_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G134gat), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n810_), .A2(G134gat), .A3(new_n624_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1343gat));
  NOR4_X1   g639(.A1(new_n630_), .A2(new_n369_), .A3(new_n410_), .A4(new_n438_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n815_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n565_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n341_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n736_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n342_), .ZN(G1345gat));
  NOR2_X1   g645(.A1(new_n842_), .A2(new_n583_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  INV_X1    g648(.A(new_n842_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n850_), .A2(G162gat), .A3(new_n669_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G162gat), .B1(new_n850_), .B2(new_n625_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  NOR3_X1   g652(.A1(new_n326_), .A2(new_n370_), .A3(new_n412_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n826_), .A2(new_n564_), .A3(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT62), .B(G169gat), .C1(new_n855_), .C2(KEYINPUT22), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n825_), .A2(new_n565_), .A3(new_n640_), .A4(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT22), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n229_), .B1(new_n859_), .B2(new_n857_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(G1348gat));
  NAND3_X1  g662(.A1(new_n815_), .A2(new_n438_), .A3(new_n854_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n736_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n230_), .ZN(G1349gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n583_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n280_), .A2(KEYINPUT123), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n220_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT123), .A2(G183gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n867_), .B2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n864_), .B2(new_n617_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n625_), .A2(new_n221_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1351gat));
  NOR2_X1   g673(.A1(new_n438_), .A2(new_n435_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n630_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n825_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n564_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n203_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n877_), .A2(new_n880_), .A3(G197gat), .A4(new_n564_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n203_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n877_), .A2(new_n527_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n205_), .A2(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT125), .B(G204gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n884_), .B2(new_n887_), .ZN(G1353gat));
  AOI21_X1  g687(.A(new_n583_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n877_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT126), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n890_), .B(new_n892_), .ZN(G1354gat));
  NAND2_X1  g692(.A1(new_n877_), .A2(new_n618_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G218gat), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n825_), .A2(G218gat), .A3(new_n624_), .A4(new_n876_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(KEYINPUT127), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n877_), .B2(new_n618_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n901_), .B2(new_n896_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n902_), .ZN(G1355gat));
endmodule


