//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT82), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n208_));
  INV_X1    g007(.A(new_n206_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT85), .Z(new_n216_));
  INV_X1    g015(.A(G141gat), .ZN(new_n217_));
  INV_X1    g016(.A(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT3), .ZN(new_n220_));
  OR3_X1    g019(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n217_), .A2(new_n218_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n220_), .B(new_n221_), .C1(new_n222_), .C2(KEYINPUT2), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n213_), .B(new_n214_), .C1(new_n216_), .C2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT84), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n225_), .A2(KEYINPUT84), .A3(new_n227_), .A4(new_n214_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n222_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n219_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n208_), .A2(new_n212_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n207_), .A2(new_n230_), .A3(new_n224_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n203_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G85gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G57gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n202_), .A3(new_n235_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n232_), .A2(new_n235_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT92), .A3(new_n202_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(new_n241_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT94), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n242_), .B(KEYINPUT92), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n250_), .A2(KEYINPUT94), .A3(new_n241_), .A4(new_n237_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n241_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n236_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n232_), .A2(new_n233_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n202_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n252_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n249_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT95), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G169gat), .ZN(new_n260_));
  INV_X1    g059(.A(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT80), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(G183gat), .B2(G190gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G169gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n261_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT24), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(G183gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT77), .Z(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n279_), .A2(KEYINPUT78), .A3(KEYINPUT26), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT26), .B1(new_n279_), .B2(KEYINPUT78), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(G183gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n275_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n268_), .B1(new_n274_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n208_), .A2(new_n212_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n288_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295_));
  INV_X1    g094(.A(G43gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G15gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n297_), .B(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n294_), .B1(new_n293_), .B2(new_n300_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n292_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n293_), .A2(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT31), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n306_), .A2(new_n301_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT95), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n249_), .A2(new_n257_), .A3(new_n309_), .A4(new_n251_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n259_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT87), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT21), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G197gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(KEYINPUT86), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n318_), .B1(new_n322_), .B2(KEYINPUT88), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n316_), .B(new_n325_), .C1(KEYINPUT88), .C2(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n285_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n277_), .A2(new_n282_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT26), .B(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n272_), .A2(new_n332_), .A3(new_n275_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT90), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n264_), .B(KEYINPUT91), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n267_), .A2(new_n262_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n329_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n314_), .B1(new_n328_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT18), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n285_), .B2(new_n327_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n314_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n334_), .A2(new_n329_), .A3(new_n336_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n338_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n329_), .A2(new_n336_), .A3(new_n333_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n328_), .A2(new_n337_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT27), .B(new_n348_), .C1(new_n352_), .C2(new_n342_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT96), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n342_), .B1(new_n338_), .B2(new_n347_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n348_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AOI211_X1 g158(.A(KEYINPUT96), .B(KEYINPUT27), .C1(new_n356_), .C2(new_n348_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n353_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT28), .Z(new_n363_));
  AOI21_X1  g162(.A(new_n329_), .B1(KEYINPUT29), .B2(new_n231_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(G78gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G106gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n365_), .B(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n361_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n311_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n259_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n374_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n379_), .B(new_n353_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT97), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n247_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n348_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n355_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n202_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n241_), .B1(new_n245_), .B2(new_n203_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n383_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n247_), .A2(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n344_), .A2(new_n349_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n314_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n351_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n314_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT93), .B1(new_n352_), .B2(new_n396_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n338_), .A2(new_n396_), .A3(new_n347_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n389_), .A2(new_n390_), .B1(new_n401_), .B2(new_n258_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n259_), .A2(new_n310_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n353_), .B(new_n374_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n402_), .A2(new_n374_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n308_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n377_), .A2(new_n381_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G120gat), .B(G148gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT5), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G176gat), .B(G204gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G85gat), .B(G92gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n419_));
  INV_X1    g218(.A(G99gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n369_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n413_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT8), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n413_), .A2(KEYINPUT9), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT9), .ZN(new_n428_));
  INV_X1    g227(.A(G85gat), .ZN(new_n429_));
  INV_X1    g228(.A(G92gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n428_), .A2(new_n431_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n432_));
  OR2_X1    g231(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n369_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n433_), .A2(KEYINPUT64), .A3(new_n369_), .A4(new_n434_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n427_), .A2(new_n432_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT8), .B(new_n413_), .C1(new_n418_), .C2(new_n423_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n426_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G78gat), .ZN(new_n442_));
  INV_X1    g241(.A(G64gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G57gat), .ZN(new_n444_));
  INV_X1    g243(.A(G57gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G64gat), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n442_), .A2(KEYINPUT11), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(KEYINPUT11), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n367_), .A2(G71gat), .ZN(new_n449_));
  INV_X1    g248(.A(G71gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G78gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT11), .B1(new_n444_), .B2(new_n446_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n447_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT12), .B1(new_n441_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n441_), .A2(new_n456_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G230gat), .A2(G233gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n447_), .B(new_n462_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n461_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT66), .B1(new_n464_), .B2(new_n441_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n463_), .A2(KEYINPUT12), .ZN(new_n466_));
  AND4_X1   g265(.A1(KEYINPUT66), .A2(new_n466_), .A3(new_n441_), .A4(new_n461_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n459_), .B(new_n460_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n460_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n426_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n455_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n471_), .B2(new_n458_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n412_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n473_), .B(KEYINPUT67), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n468_), .A2(new_n472_), .A3(new_n412_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT68), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT74), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT74), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G15gat), .A2(G22gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G15gat), .A2(G22gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(G1gat), .B2(G8gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT73), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n495_), .B1(new_n502_), .B2(new_n491_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G1gat), .B(G8gat), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n494_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT74), .B1(new_n492_), .B2(new_n493_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n495_), .A3(new_n491_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT70), .ZN(new_n513_));
  INV_X1    g312(.A(G36gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G29gat), .ZN(new_n515_));
  INV_X1    g314(.A(G29gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G36gat), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n515_), .A2(new_n517_), .A3(KEYINPUT70), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n511_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n517_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(KEYINPUT70), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n510_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n506_), .A2(new_n509_), .A3(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n505_), .B1(new_n494_), .B2(new_n503_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n507_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n485_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(KEYINPUT15), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n534_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n528_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n484_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT75), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n531_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(KEYINPUT76), .A3(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n407_), .A2(new_n483_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n532_), .A2(new_n441_), .A3(new_n534_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n470_), .A2(new_n525_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(new_n560_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n554_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n566_), .A2(KEYINPUT72), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT72), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n564_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .A4(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(KEYINPUT37), .C1(new_n571_), .C2(new_n566_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n566_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT71), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n528_), .A2(new_n529_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n455_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(KEYINPUT65), .A3(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(KEYINPUT17), .B2(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n582_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n578_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n550_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n488_), .A3(new_n403_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT38), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n567_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n593_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n550_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n403_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(G1324gat));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n489_), .A3(new_n361_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  INV_X1    g407(.A(new_n603_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n361_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n610_), .B2(G8gat), .ZN(new_n611_));
  AOI211_X1 g410(.A(KEYINPUT39), .B(new_n489_), .C1(new_n609_), .C2(new_n361_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n607_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(KEYINPUT40), .B(new_n607_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n596_), .A2(new_n618_), .A3(new_n308_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT98), .Z(new_n620_));
  OAI21_X1  g419(.A(G15gat), .B1(new_n603_), .B2(new_n406_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT41), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n603_), .B2(new_n379_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n596_), .A2(new_n626_), .A3(new_n374_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(G1327gat));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n407_), .B2(new_n578_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n377_), .A2(new_n381_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n405_), .A2(new_n406_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(KEYINPUT44), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n483_), .A2(new_n549_), .A3(new_n593_), .A4(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n637_), .A3(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(KEYINPUT44), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(new_n639_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n516_), .B1(new_n644_), .B2(new_n403_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n599_), .A2(new_n593_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n550_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n403_), .A2(new_n516_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT100), .Z(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT101), .B1(new_n645_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n604_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n654_));
  OAI221_X1 g453(.A(new_n653_), .B1(new_n648_), .B2(new_n650_), .C1(new_n654_), .C2(new_n516_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n514_), .B1(new_n644_), .B2(new_n361_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n361_), .B(KEYINPUT102), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n647_), .A2(new_n514_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n359_), .A2(new_n360_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n641_), .A2(new_n643_), .B1(new_n666_), .B2(new_n353_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n665_), .B(KEYINPUT46), .C1(new_n667_), .C2(new_n514_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(G1329gat));
  AOI21_X1  g468(.A(G43gat), .B1(new_n647_), .B2(new_n308_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n406_), .A2(new_n296_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n644_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n647_), .B2(new_n374_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n374_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n644_), .B2(new_n676_), .ZN(G1331gat));
  AND2_X1   g476(.A1(new_n547_), .A2(new_n548_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n407_), .A2(new_n482_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n595_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT103), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n604_), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n602_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n604_), .A2(new_n445_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1332gat));
  NAND3_X1  g489(.A1(new_n681_), .A2(new_n443_), .A3(new_n660_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT48), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n660_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G64gat), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT48), .B(new_n443_), .C1(new_n688_), .C2(new_n660_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1333gat));
  NAND3_X1  g495(.A1(new_n681_), .A2(new_n450_), .A3(new_n308_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n688_), .A2(new_n308_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT49), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(G71gat), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G71gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1334gat));
  NAND3_X1  g501(.A1(new_n681_), .A2(new_n367_), .A3(new_n374_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n688_), .A2(new_n374_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G78gat), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT50), .B(new_n367_), .C1(new_n688_), .C2(new_n374_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1335gat));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n636_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n629_), .A2(new_n635_), .A3(KEYINPUT106), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n482_), .A2(new_n678_), .A3(new_n593_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n604_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n679_), .A2(new_n646_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n429_), .A3(new_n403_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n713_), .B2(new_n659_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n430_), .A3(new_n361_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1337gat));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n710_), .A2(new_n308_), .A3(new_n711_), .A4(new_n712_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G99gat), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n715_), .A2(new_n433_), .A3(new_n434_), .A4(new_n308_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n722_), .B(new_n723_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  AND4_X1   g526(.A1(new_n721_), .A2(new_n725_), .A3(KEYINPUT51), .A4(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n715_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n712_), .A2(new_n374_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n369_), .B1(new_n732_), .B2(KEYINPUT108), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734_));
  INV_X1    g533(.A(new_n731_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n407_), .A2(KEYINPUT43), .A3(new_n578_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n633_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n733_), .A2(new_n734_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n734_), .B1(new_n733_), .B2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n730_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n730_), .B(new_n744_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1339gat));
  NOR2_X1   g547(.A1(new_n594_), .A2(new_n678_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n482_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n750_), .B(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n484_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n535_), .A2(new_n485_), .A3(new_n536_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n543_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n476_), .A2(new_n546_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n468_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n459_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT66), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n461_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n470_), .B2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n466_), .A2(new_n441_), .A3(KEYINPUT66), .A4(new_n461_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT113), .A3(new_n459_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n469_), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n468_), .A2(KEYINPUT112), .A3(new_n759_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n770_), .A2(KEYINPUT55), .A3(new_n460_), .A4(new_n459_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT114), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n411_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT56), .B(new_n411_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n758_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n754_), .B(new_n634_), .C1(new_n781_), .C2(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n758_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n780_), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n458_), .B(new_n457_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n787_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n460_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n775_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(new_n772_), .A3(new_n762_), .A4(new_n773_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n411_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n754_), .B1(new_n796_), .B2(new_n634_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT117), .B1(new_n784_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n634_), .B1(new_n781_), .B2(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n757_), .A2(new_n546_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n678_), .A2(new_n805_), .A3(new_n476_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT68), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n475_), .B(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n808_), .B2(new_n549_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n779_), .A2(new_n780_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n812_), .A2(new_n600_), .B1(new_n813_), .B2(KEYINPUT57), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n806_), .A2(new_n809_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n599_), .B(new_n815_), .C1(new_n817_), .C2(new_n804_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n798_), .A2(new_n802_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n753_), .B1(new_n820_), .B2(new_n601_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n604_), .A2(new_n406_), .A3(new_n380_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n800_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n593_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(new_n822_), .C1(new_n827_), .C2(new_n753_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n678_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G113gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n820_), .A2(new_n601_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n753_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n823_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n549_), .A2(G113gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n830_), .B1(new_n834_), .B2(new_n835_), .ZN(G1340gat));
  OAI211_X1 g635(.A(new_n483_), .B(new_n828_), .C1(new_n833_), .C2(new_n825_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n482_), .B2(G120gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n824_), .A2(KEYINPUT118), .A3(new_n483_), .A4(new_n828_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G120gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n833_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1341gat));
  NAND3_X1  g646(.A1(new_n824_), .A2(new_n593_), .A3(new_n828_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G127gat), .ZN(new_n849_));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n833_), .A2(new_n850_), .A3(new_n593_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n849_), .A2(KEYINPUT119), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1342gat));
  NAND3_X1  g655(.A1(new_n824_), .A2(new_n634_), .A3(new_n828_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G134gat), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n599_), .A2(G134gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n834_), .B2(new_n859_), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n308_), .A2(new_n379_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n660_), .A2(new_n604_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n821_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n678_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(KEYINPUT121), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(G141gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n867_), .A2(new_n868_), .A3(new_n870_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n865_), .A2(new_n483_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n865_), .A2(new_n593_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n865_), .A2(KEYINPUT122), .A3(new_n593_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(new_n865_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n884_), .A2(G162gat), .A3(new_n599_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G162gat), .B1(new_n884_), .B2(new_n578_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n827_), .A2(new_n753_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n660_), .A2(KEYINPUT123), .A3(new_n311_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n659_), .B2(new_n378_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n374_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(new_n678_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n888_), .B1(new_n895_), .B2(new_n269_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n260_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT124), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n896_), .A2(new_n898_), .A3(new_n901_), .A4(new_n897_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1348gat));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n826_), .A2(KEYINPUT117), .B1(new_n814_), .B2(new_n818_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n593_), .B1(new_n905_), .B2(new_n802_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n904_), .B(new_n379_), .C1(new_n906_), .C2(new_n753_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT125), .B1(new_n821_), .B2(new_n374_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n890_), .A2(new_n892_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n482_), .A2(new_n261_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .A4(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n889_), .A2(new_n893_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n261_), .B1(new_n912_), .B2(new_n482_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1349gat));
  AND4_X1   g713(.A1(new_n593_), .A2(new_n907_), .A3(new_n908_), .A4(new_n909_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G183gat), .B1(new_n915_), .B2(KEYINPUT126), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n601_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n912_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n601_), .A2(new_n330_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n916_), .A2(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n912_), .B2(new_n578_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n600_), .A2(new_n331_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n912_), .B2(new_n924_), .ZN(G1351gat));
  NAND3_X1  g724(.A1(new_n660_), .A2(new_n604_), .A3(new_n861_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n821_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n678_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n483_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g730(.A(new_n601_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n927_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT127), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n927_), .A2(new_n935_), .A3(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(new_n927_), .ZN(new_n940_));
  OR3_X1    g739(.A1(new_n940_), .A2(G218gat), .A3(new_n599_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G218gat), .B1(new_n940_), .B2(new_n578_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1355gat));
endmodule


