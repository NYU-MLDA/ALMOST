//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(G22gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G1gat), .B(G8gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT79), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n209_), .A2(new_n212_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n209_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n221_), .A2(new_n213_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT80), .B1(new_n227_), .B2(KEYINPUT81), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n232_), .B2(new_n227_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT12), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n235_), .A2(KEYINPUT69), .ZN(new_n236_));
  XOR2_X1   g035(.A(G85gat), .B(G92gat), .Z(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(KEYINPUT9), .A2(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(G92gat), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT9), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244_));
  AND3_X1   g043(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT65), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n243_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT7), .ZN(new_n256_));
  INV_X1    g055(.A(G99gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n239_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n245_), .A2(new_n246_), .A3(new_n244_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT65), .B1(new_n250_), .B2(new_n251_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT8), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n237_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT66), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n260_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n266_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n258_), .A2(new_n250_), .A3(new_n251_), .A4(new_n259_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n265_), .B1(new_n273_), .B2(new_n237_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT67), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n255_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(G57gat), .A2(G64gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G57gat), .A2(G64gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n280_));
  INV_X1    g079(.A(G71gat), .ZN(new_n281_));
  INV_X1    g080(.A(G78gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n279_), .A2(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT68), .B1(new_n279_), .B2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G71gat), .A2(G78gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(KEYINPUT11), .C1(new_n277_), .C2(new_n278_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n282_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n285_), .B(new_n289_), .C1(new_n290_), .C2(KEYINPUT11), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n290_), .B2(KEYINPUT11), .ZN(new_n292_));
  INV_X1    g091(.A(new_n287_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n288_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n236_), .B1(new_n276_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT64), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n235_), .A2(KEYINPUT69), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n273_), .A2(new_n237_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT8), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT67), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n264_), .A2(KEYINPUT66), .A3(new_n267_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n270_), .B1(new_n269_), .B2(new_n266_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(KEYINPUT8), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n254_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n295_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n300_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n299_), .B(new_n295_), .C1(new_n308_), .C2(new_n254_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n296_), .B(new_n298_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n276_), .A2(new_n295_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n310_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n313_), .B1(new_n298_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G204gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT5), .B(G176gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT70), .Z(new_n322_));
  AND2_X1   g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n317_), .A2(new_n321_), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT13), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT13), .B1(new_n323_), .B2(new_n324_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n234_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G231gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n209_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(new_n295_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT77), .Z(new_n332_));
  XNOR2_X1  g131(.A(G127gat), .B(G155gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G211gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT16), .B(G183gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT17), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT78), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT17), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n331_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n328_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n346_));
  OAI21_X1  g145(.A(G169gat), .B1(new_n346_), .B2(G176gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT22), .B(G169gat), .Z(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT85), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n353_));
  AND2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(new_n354_), .ZN(new_n357_));
  MUX2_X1   g156(.A(new_n355_), .B(new_n357_), .S(KEYINPUT86), .Z(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(G183gat), .B2(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n356_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT83), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(KEYINPUT83), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(new_n354_), .C2(new_n353_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT25), .B(G183gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n366_), .A2(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT24), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n364_), .B(new_n370_), .C1(new_n369_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n360_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(G197gat), .B(G204gat), .Z(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(KEYINPUT21), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(KEYINPUT21), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n360_), .A2(KEYINPUT87), .A3(new_n373_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n372_), .B(KEYINPUT93), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n358_), .B(new_n370_), .C1(new_n369_), .C2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n364_), .B1(G183gat), .B2(G190gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT96), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT94), .A2(G169gat), .A3(G176gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n349_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT95), .Z(new_n392_));
  OAI21_X1  g191(.A(new_n385_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n381_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT19), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT97), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n376_), .A2(new_n382_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n394_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n398_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n393_), .A2(new_n394_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(KEYINPUT97), .A3(new_n398_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT18), .B(G64gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n401_), .A2(new_n406_), .A3(new_n407_), .A4(new_n412_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT27), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT100), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G155gat), .B(G162gat), .Z(new_n419_));
  NAND2_X1  g218(.A1(G141gat), .A2(G148gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT2), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(KEYINPUT90), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(KEYINPUT90), .ZN(new_n423_));
  MUX2_X1   g222(.A(new_n420_), .B(new_n422_), .S(new_n423_), .Z(new_n424_));
  OR2_X1    g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT3), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n419_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n419_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n420_), .A3(new_n425_), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(KEYINPUT29), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT28), .B(G22gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G50gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n433_), .B(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT91), .B1(G228gat), .B2(G233gat), .ZN(new_n437_));
  AND3_X1   g236(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n437_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n381_), .B1(new_n432_), .B2(KEYINPUT29), .ZN(new_n440_));
  MUX2_X1   g239(.A(new_n437_), .B(new_n439_), .S(new_n440_), .Z(new_n441_));
  XOR2_X1   g240(.A(G78gat), .B(G106gat), .Z(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n443_), .B2(KEYINPUT92), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n441_), .B(new_n442_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G120gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(G127gat), .B(G134gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT89), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n402_), .A2(KEYINPUT30), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n402_), .A2(KEYINPUT30), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n456_), .A2(G71gat), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n402_), .A2(KEYINPUT30), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n281_), .B1(new_n459_), .B2(new_n455_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n454_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(G71gat), .B1(new_n456_), .B2(new_n457_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n454_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n281_), .A3(new_n455_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT88), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G99gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n447_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n461_), .A2(new_n465_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n446_), .A3(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n432_), .B(new_n450_), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT4), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n432_), .A2(new_n450_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(KEYINPUT4), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(new_n241_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n396_), .A2(new_n398_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n405_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n404_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n413_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT27), .A3(new_n415_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n418_), .A2(new_n477_), .A3(new_n494_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT98), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n408_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n501_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n497_), .A2(KEYINPUT99), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT99), .B1(new_n497_), .B2(new_n504_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n503_), .B(new_n493_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n492_), .B(KEYINPUT33), .ZN(new_n508_));
  INV_X1    g307(.A(new_n482_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n478_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n489_), .B(new_n510_), .C1(new_n481_), .C2(new_n509_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n414_), .A2(new_n508_), .A3(new_n415_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n475_), .A2(new_n469_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n446_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n345_), .B1(new_n500_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n276_), .A2(new_n212_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n309_), .A2(new_n220_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT34), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n517_), .B(new_n518_), .C1(KEYINPUT35), .C2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  INV_X1    g323(.A(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT71), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n521_), .A2(new_n522_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT72), .B1(new_n533_), .B2(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT37), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(KEYINPUT73), .A3(new_n534_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n532_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n539_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n516_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n493_), .B(KEYINPUT101), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n204_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT103), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n542_), .A2(new_n532_), .A3(new_n543_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n516_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n204_), .B1(new_n557_), .B2(new_n493_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(KEYINPUT103), .A3(new_n554_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n559_), .B(new_n560_), .C1(new_n554_), .C2(new_n552_), .ZN(G1324gat));
  INV_X1    g360(.A(KEYINPUT40), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n418_), .A2(new_n499_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n550_), .A2(new_n205_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT104), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n205_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT39), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT40), .A3(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(G1325gat));
  INV_X1    g371(.A(G15gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n514_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n557_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT41), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n550_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1326gat));
  INV_X1    g377(.A(G22gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n550_), .A2(new_n579_), .A3(new_n447_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n557_), .B2(new_n447_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT105), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT42), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n582_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n580_), .B1(new_n586_), .B2(new_n587_), .ZN(G1327gat));
  NOR2_X1   g387(.A1(new_n416_), .A2(new_n417_), .ZN(new_n589_));
  AOI211_X1 g388(.A(KEYINPUT100), .B(KEYINPUT27), .C1(new_n414_), .C2(new_n415_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n494_), .B(new_n499_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n470_), .A2(new_n447_), .A3(new_n471_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n446_), .B1(new_n475_), .B2(new_n469_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n515_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT43), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n548_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n595_), .B2(new_n548_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n328_), .B(new_n343_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT44), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n548_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT43), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n596_), .A3(new_n548_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT44), .A3(new_n328_), .A4(new_n343_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n606_), .A3(new_n551_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G29gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n556_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n595_), .A2(new_n609_), .A3(new_n328_), .A4(new_n343_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n494_), .A2(G29gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT106), .Z(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n610_), .B2(new_n612_), .ZN(G1328gat));
  INV_X1    g412(.A(KEYINPUT107), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(G36gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n563_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT45), .ZN(new_n617_));
  INV_X1    g416(.A(new_n563_), .ZN(new_n618_));
  NOR4_X1   g417(.A1(new_n610_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n616_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n556_), .B1(new_n500_), .B2(new_n515_), .ZN(new_n621_));
  INV_X1    g420(.A(G36gat), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n328_), .A4(new_n343_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT107), .B1(new_n623_), .B2(new_n618_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n614_), .A3(new_n563_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT45), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n601_), .A2(new_n606_), .A3(new_n563_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G36gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT108), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT46), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n627_), .A2(new_n629_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n631_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n617_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n624_), .A2(new_n625_), .A3(KEYINPUT45), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n618_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n622_), .B1(new_n638_), .B2(new_n606_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n633_), .B(new_n634_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n632_), .A2(new_n640_), .ZN(G1329gat));
  NAND4_X1  g440(.A1(new_n601_), .A2(new_n606_), .A3(G43gat), .A4(new_n574_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n610_), .A2(new_n514_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(G43gat), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g444(.A1(new_n610_), .A2(new_n446_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(G50gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n606_), .A2(G50gat), .A3(new_n447_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n649_), .B2(new_n601_), .ZN(G1331gat));
  AOI21_X1  g449(.A(new_n343_), .B1(new_n500_), .B2(new_n515_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n327_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n233_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n651_), .A2(new_n549_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G57gat), .B1(new_n654_), .B2(new_n551_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n556_), .A3(new_n653_), .ZN(new_n656_));
  INV_X1    g455(.A(G57gat), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n494_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1332gat));
  OAI21_X1  g458(.A(G64gat), .B1(new_n656_), .B2(new_n618_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT48), .ZN(new_n661_));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n654_), .A2(new_n662_), .A3(new_n563_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1333gat));
  OAI21_X1  g463(.A(G71gat), .B1(new_n656_), .B2(new_n514_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT49), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n654_), .A2(new_n281_), .A3(new_n574_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1334gat));
  OAI21_X1  g467(.A(G78gat), .B1(new_n656_), .B2(new_n446_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n654_), .A2(new_n282_), .A3(new_n447_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1335gat));
  NAND2_X1  g472(.A1(new_n653_), .A2(new_n343_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n621_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G85gat), .B1(new_n676_), .B2(new_n551_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n605_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n603_), .A2(KEYINPUT110), .A3(new_n604_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n675_), .A3(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n494_), .A2(new_n241_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n677_), .B1(new_n681_), .B2(new_n682_), .ZN(G1336gat));
  NAND4_X1  g482(.A1(new_n679_), .A2(new_n563_), .A3(new_n675_), .A4(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G92gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n676_), .A2(new_n242_), .A3(new_n563_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT111), .ZN(G1337gat));
  NAND4_X1  g487(.A1(new_n679_), .A2(new_n574_), .A3(new_n675_), .A4(new_n680_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G99gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n238_), .A3(new_n574_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g492(.A1(new_n652_), .A2(new_n233_), .A3(new_n446_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n621_), .A2(new_n239_), .A3(new_n343_), .A4(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n605_), .A2(new_n343_), .A3(new_n694_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT52), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G106gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G106gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g500(.A1(new_n618_), .A2(new_n551_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n476_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n327_), .A2(new_n343_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n234_), .B(new_n706_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT54), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n707_), .A2(KEYINPUT54), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n313_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n315_), .A2(new_n299_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n309_), .A2(new_n310_), .A3(new_n300_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT55), .A3(new_n298_), .A4(new_n296_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n296_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n298_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n313_), .A2(KEYINPUT113), .A3(new_n714_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n717_), .A2(new_n721_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT114), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n721_), .A2(new_n724_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n717_), .A4(new_n725_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n322_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT115), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n324_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n735_), .A2(new_n233_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n216_), .A2(new_n217_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n227_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n227_), .B2(new_n224_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n323_), .A2(new_n324_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n609_), .B1(new_n738_), .B2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT57), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n737_), .A2(new_n233_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n324_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n609_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n747_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n732_), .A2(new_n734_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(KEYINPUT118), .A3(new_n734_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n313_), .A2(KEYINPUT113), .A3(new_n714_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT113), .B1(new_n313_), .B2(new_n714_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n730_), .B1(new_n760_), .B2(new_n729_), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n728_), .A2(new_n758_), .A3(new_n759_), .A4(KEYINPUT114), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n322_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n756_), .A2(new_n757_), .A3(new_n764_), .A4(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n742_), .A2(new_n324_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(KEYINPUT58), .A3(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n548_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n344_), .B1(new_n753_), .B2(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n704_), .B(new_n705_), .C1(new_n713_), .C2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n702_), .A2(new_n476_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n746_), .B2(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n751_), .B1(new_n750_), .B2(new_n609_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n738_), .A2(new_n745_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n556_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n778_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n343_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n777_), .B1(new_n785_), .B2(new_n712_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n775_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT120), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n775_), .B(new_n790_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n789_), .A2(G113gat), .A3(new_n233_), .A4(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(G113gat), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n767_), .A2(KEYINPUT58), .A3(new_n768_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT58), .B1(new_n767_), .B2(new_n768_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n796_), .A2(new_n548_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n747_), .B2(new_n752_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n344_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n776_), .B1(new_n799_), .B2(new_n713_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n793_), .B1(new_n800_), .B2(new_n234_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n792_), .A2(new_n801_), .ZN(G1340gat));
  INV_X1    g601(.A(KEYINPUT60), .ZN(new_n803_));
  AOI21_X1  g602(.A(G120gat), .B1(new_n327_), .B2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n803_), .A2(G120gat), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n800_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT121), .ZN(new_n807_));
  OAI21_X1  g606(.A(G120gat), .B1(new_n788_), .B2(new_n652_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1341gat));
  NAND4_X1  g608(.A1(new_n789_), .A2(G127gat), .A3(new_n344_), .A4(new_n791_), .ZN(new_n810_));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n800_), .B2(new_n343_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1342gat));
  NAND4_X1  g612(.A1(new_n789_), .A2(G134gat), .A3(new_n548_), .A4(new_n791_), .ZN(new_n814_));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n800_), .B2(new_n556_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1343gat));
  NAND3_X1  g616(.A1(new_n618_), .A2(new_n551_), .A3(new_n593_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n785_), .B2(new_n712_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n233_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT122), .B(G141gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1344gat));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n327_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n344_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  NAND2_X1  g626(.A1(new_n548_), .A2(G162gat), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT124), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n819_), .A2(new_n829_), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT123), .B(G162gat), .C1(new_n819_), .C2(new_n609_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n832_));
  INV_X1    g631(.A(new_n818_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n609_), .B(new_n833_), .C1(new_n799_), .C2(new_n713_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n525_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n830_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT125), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n830_), .C1(new_n831_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1347gat));
  INV_X1    g639(.A(G169gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n713_), .A2(new_n774_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n618_), .A2(new_n551_), .A3(new_n476_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n844_), .B2(new_n233_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n842_), .A2(new_n234_), .A3(new_n348_), .A4(new_n843_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT62), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(KEYINPUT62), .B2(new_n845_), .ZN(G1348gat));
  AOI21_X1  g647(.A(G176gat), .B1(new_n844_), .B2(new_n327_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n785_), .B2(new_n712_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n327_), .A2(G176gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  AOI21_X1  g651(.A(G183gat), .B1(new_n850_), .B2(new_n344_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n343_), .A2(new_n366_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n844_), .B2(new_n854_), .ZN(G1350gat));
  NAND3_X1  g654(.A1(new_n844_), .A2(new_n609_), .A3(new_n367_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n842_), .A2(new_n549_), .A3(new_n843_), .ZN(new_n857_));
  INV_X1    g656(.A(G190gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1351gat));
  NAND2_X1  g658(.A1(new_n593_), .A2(new_n494_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT126), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(KEYINPUT126), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n563_), .A2(new_n862_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n861_), .B(new_n863_), .C1(new_n785_), .C2(new_n712_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n233_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n327_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n344_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  AND2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n869_), .B2(new_n870_), .ZN(G1354gat));
  AOI21_X1  g672(.A(G218gat), .B1(new_n864_), .B2(new_n609_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n548_), .A2(G218gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT127), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n864_), .B2(new_n876_), .ZN(G1355gat));
endmodule


