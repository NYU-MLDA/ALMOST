//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n986_, new_n987_, new_n988_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1001_, new_n1002_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT91), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n206_), .B2(new_n205_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT86), .B1(new_n216_), .B2(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G190gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(G183gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT86), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n215_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT87), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(new_n215_), .C1(new_n222_), .C2(new_n226_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(G183gat), .A3(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT88), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(new_n232_), .A3(G183gat), .A4(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n223_), .B2(new_n218_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n231_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n230_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n233_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n245_));
  NOR3_X1   g044(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G15gat), .B(G43gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT90), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n252_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G71gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n255_), .A2(new_n257_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n210_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n209_), .A3(new_n258_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  OR3_X1    g063(.A1(KEYINPUT94), .A2(G155gat), .A3(G162gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT94), .B1(G155gat), .B2(G162gat), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n265_), .A2(new_n266_), .B1(G155gat), .B2(G162gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  INV_X1    g067(.A(G141gat), .ZN(new_n269_));
  INV_X1    g068(.A(G148gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .A4(KEYINPUT95), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT95), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n273_), .A2(G141gat), .A3(G148gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n271_), .B(new_n272_), .C1(new_n274_), .C2(new_n268_), .ZN(new_n275_));
  AND3_X1   g074(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT92), .B1(G141gat), .B2(G148gat), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT2), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n267_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n266_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(KEYINPUT94), .A2(G155gat), .A3(G162gat), .ZN(new_n281_));
  AND3_X1   g080(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n280_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n276_), .A2(new_n277_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(new_n205_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT100), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n205_), .B1(new_n279_), .B2(new_n289_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n279_), .A2(new_n289_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n205_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT100), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT4), .B1(new_n293_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT101), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(new_n295_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(KEYINPUT4), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(KEYINPUT100), .A3(new_n290_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n306_), .B2(new_n297_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n305_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n297_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n303_), .B1(new_n315_), .B2(KEYINPUT4), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(new_n307_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n317_), .B2(new_n311_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G78gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G106gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G22gat), .B(G50gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n279_), .A2(new_n289_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT28), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT97), .B1(new_n333_), .B2(G197gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT97), .ZN(new_n335_));
  INV_X1    g134(.A(G197gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(G204gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(G197gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n332_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT96), .B1(new_n333_), .B2(G197gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT96), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n336_), .A3(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n343_), .A3(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT21), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n334_), .A2(new_n337_), .A3(new_n331_), .A4(new_n338_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n330_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n340_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n329_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n329_), .B2(new_n353_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n325_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n354_), .A3(new_n324_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n241_), .B1(KEYINPUT24), .B2(new_n213_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT25), .B(G183gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n215_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(KEYINPUT98), .A3(new_n215_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n242_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n245_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT99), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n379_), .A2(new_n246_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT99), .B1(new_n247_), .B2(new_n245_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT104), .ZN(new_n385_));
  INV_X1    g184(.A(new_n348_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n386_), .A2(new_n345_), .B1(new_n339_), .B2(new_n332_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT104), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n249_), .B2(new_n349_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n368_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n349_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n240_), .A2(new_n387_), .A3(new_n248_), .ZN(new_n395_));
  AND4_X1   g194(.A1(KEYINPUT20), .A2(new_n394_), .A3(new_n368_), .A4(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n365_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n365_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n387_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n367_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT20), .A4(new_n367_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n398_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n397_), .A2(KEYINPUT27), .A3(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n377_), .A2(new_n383_), .A3(new_n349_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n387_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n391_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n401_), .B(new_n365_), .C1(new_n407_), .C2(new_n367_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT27), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n404_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n264_), .A2(new_n319_), .A3(new_n361_), .A4(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n360_), .B(new_n314_), .C1(new_n311_), .C2(new_n317_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n404_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n301_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n293_), .B2(new_n298_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n311_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT33), .B1(new_n417_), .B2(new_n316_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n305_), .A2(new_n313_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n301_), .B1(new_n293_), .B2(new_n298_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n312_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n415_), .B1(new_n302_), .B2(KEYINPUT4), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n315_), .B2(KEYINPUT4), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT102), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n299_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT102), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n311_), .B1(new_n315_), .B2(new_n301_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n409_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT103), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n409_), .A2(new_n421_), .A3(new_n432_), .A4(KEYINPUT103), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n393_), .A2(new_n396_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n318_), .B(new_n438_), .C1(new_n439_), .C2(new_n437_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n414_), .B1(new_n441_), .B2(new_n361_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n412_), .B1(new_n442_), .B2(new_n264_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G230gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G64gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G78gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n449_));
  XOR2_X1   g248(.A(G71gat), .B(G78gat), .Z(new_n450_));
  INV_X1    g249(.A(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G57gat), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G64gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT11), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n446_), .B(new_n449_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n452_), .A2(new_n454_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n455_), .A3(new_n450_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n446_), .B1(new_n463_), .B2(new_n449_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467_));
  INV_X1    g266(.A(G85gat), .ZN(new_n468_));
  INV_X1    g267(.A(G92gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n467_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n479_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n466_), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n466_), .B1(new_n486_), .B2(new_n472_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT65), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n479_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n487_), .B1(KEYINPUT66), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n489_), .A2(new_n495_), .A3(new_n479_), .A4(new_n492_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n485_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n489_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n470_), .B1(new_n503_), .B2(new_n471_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n471_), .A2(new_n503_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n471_), .A2(KEYINPUT64), .A3(new_n503_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n502_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(KEYINPUT69), .B(new_n465_), .C1(new_n497_), .C2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT69), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n493_), .A2(KEYINPUT66), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT8), .B1(new_n473_), .B2(new_n474_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n496_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n475_), .A2(new_n484_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n510_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n465_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n497_), .A2(new_n510_), .A3(new_n465_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n445_), .B(new_n511_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n463_), .A2(new_n449_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT12), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n492_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT65), .B1(new_n490_), .B2(new_n491_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n507_), .A2(new_n508_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n504_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n531_), .A2(new_n534_), .A3(new_n535_), .A4(new_n501_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT70), .B1(new_n502_), .B2(new_n509_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n497_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n518_), .A2(new_n519_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n524_), .A2(new_n444_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G120gat), .B(G148gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G176gat), .B(G204gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n522_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n522_), .A2(new_n541_), .A3(KEYINPUT71), .A4(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n522_), .A2(new_n541_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n551_), .A2(new_n553_), .B1(new_n556_), .B2(new_n554_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G1gat), .B(G8gat), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G1gat), .A2(G8gat), .ZN(new_n561_));
  OR2_X1    g360(.A1(G15gat), .A2(G22gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G15gat), .A2(G22gat), .ZN(new_n563_));
  AOI221_X4 g362(.A(KEYINPUT78), .B1(new_n561_), .B2(KEYINPUT14), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G15gat), .B(G22gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(KEYINPUT14), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n564_), .A2(new_n568_), .A3(KEYINPUT79), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT79), .ZN(new_n570_));
  AND2_X1   g369(.A1(G15gat), .A2(G22gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(G15gat), .A2(G22gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n561_), .A2(KEYINPUT14), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT78), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n570_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n560_), .B1(new_n569_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT79), .B1(new_n564_), .B2(new_n568_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n559_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G29gat), .B(G36gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G43gat), .B(G50gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT83), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT83), .ZN(new_n591_));
  INV_X1    g390(.A(new_n586_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n579_), .A2(new_n559_), .A3(new_n580_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n559_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n591_), .B1(new_n595_), .B2(KEYINPUT82), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n587_), .B1(new_n590_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT83), .B1(new_n588_), .B2(new_n589_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(KEYINPUT82), .A3(new_n591_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n583_), .A4(new_n586_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n586_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n583_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT84), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n603_), .A2(new_n608_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n558_), .A2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n582_), .A2(KEYINPUT80), .ZN(new_n620_));
  AND2_X1   g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n582_), .A2(KEYINPUT80), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n525_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n526_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n627_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n625_), .A2(new_n465_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n519_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n632_), .B(KEYINPUT17), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G232gat), .A2(G233gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT34), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT35), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n518_), .A2(new_n592_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n515_), .A2(new_n517_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n536_), .A2(new_n537_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n605_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n646_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n606_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n646_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n648_), .A4(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT76), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G190gat), .B(G218gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT75), .ZN(new_n660_));
  XOR2_X1   g459(.A(G134gat), .B(G162gat), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT36), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n664_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n653_), .A2(KEYINPUT76), .A3(new_n657_), .A4(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n653_), .A2(new_n657_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n662_), .A2(new_n663_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n641_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n443_), .A2(new_n619_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n202_), .B1(new_n676_), .B2(new_n318_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT85), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n603_), .A2(new_n608_), .A3(new_n615_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n615_), .B1(new_n603_), .B2(new_n608_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n614_), .A2(KEYINPUT85), .A3(new_n616_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n443_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT73), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n558_), .B(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT77), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n672_), .A2(new_n687_), .A3(KEYINPUT37), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT37), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n665_), .A2(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(KEYINPUT77), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n691_), .A3(new_n640_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n686_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n684_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n693_), .A3(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n202_), .A3(new_n318_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n677_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n698_), .A2(new_n202_), .A3(new_n702_), .A4(new_n318_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT107), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT107), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1324gat));
  NOR2_X1   g505(.A1(new_n411_), .A2(G8gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n695_), .A2(new_n697_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G8gat), .B1(new_n674_), .B2(new_n411_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT39), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT39), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT110), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n708_), .B(new_n714_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(G1325gat));
  INV_X1    g517(.A(new_n264_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n694_), .A2(G15gat), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n676_), .A2(new_n264_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT41), .B1(new_n721_), .B2(G15gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1326gat));
  OR3_X1    g523(.A1(new_n694_), .A2(G22gat), .A3(new_n361_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n676_), .A2(new_n360_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(G22gat), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G22gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT112), .ZN(G1327gat));
  INV_X1    g530(.A(new_n558_), .ZN(new_n732_));
  AND4_X1   g531(.A1(new_n684_), .A2(new_n732_), .A3(new_n672_), .A4(new_n641_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G29gat), .B1(new_n733_), .B2(new_n318_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n688_), .A2(new_n691_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n443_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n443_), .A2(KEYINPUT113), .A3(new_n735_), .A4(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n443_), .A2(new_n736_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT43), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n619_), .A2(new_n641_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n743_), .A2(KEYINPUT44), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n745_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT44), .B1(new_n747_), .B2(KEYINPUT114), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n743_), .A2(new_n749_), .A3(new_n745_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n746_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n318_), .A2(G29gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n734_), .B1(new_n751_), .B2(new_n752_), .ZN(G1328gat));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n754_));
  INV_X1    g553(.A(G36gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n747_), .A2(KEYINPUT114), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n750_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n746_), .A2(new_n411_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n411_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n733_), .A2(new_n755_), .A3(new_n761_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT45), .Z(new_n763_));
  OAI21_X1  g562(.A(new_n754_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n762_), .B(KEYINPUT45), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n747_), .B2(new_n757_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n750_), .B2(new_n748_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT46), .B(new_n765_), .C1(new_n767_), .C2(new_n755_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n768_), .ZN(G1329gat));
  INV_X1    g568(.A(G43gat), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n719_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n772_), .B(new_n746_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n733_), .A2(new_n264_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n770_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT47), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n751_), .A2(new_n771_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1330gat));
  AOI21_X1  g580(.A(G50gat), .B1(new_n733_), .B2(new_n360_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n360_), .A2(G50gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n751_), .B2(new_n783_), .ZN(G1331gat));
  INV_X1    g583(.A(new_n686_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n683_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n443_), .A2(new_n673_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n788_), .A2(new_n453_), .A3(new_n319_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n443_), .A2(new_n618_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n732_), .A2(new_n692_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n793_), .A2(KEYINPUT115), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT115), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n318_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n789_), .B1(new_n796_), .B2(new_n453_), .ZN(G1332gat));
  OAI21_X1  g596(.A(G64gat), .B1(new_n788_), .B2(new_n411_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT48), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n793_), .A2(new_n451_), .A3(new_n761_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1333gat));
  OR3_X1    g600(.A1(new_n792_), .A2(G71gat), .A3(new_n719_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n786_), .A2(new_n264_), .A3(new_n787_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(G71gat), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(G71gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT117), .Z(G1334gat));
  OAI21_X1  g607(.A(G78gat), .B1(new_n788_), .B2(new_n361_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n361_), .A2(G78gat), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT119), .Z(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n792_), .B2(new_n813_), .ZN(G1335gat));
  NOR3_X1   g613(.A1(new_n732_), .A2(new_n617_), .A3(new_n640_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n743_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816_), .B2(new_n319_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n785_), .A2(new_n690_), .A3(new_n640_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n790_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n468_), .A3(new_n318_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(G1336gat));
  OAI21_X1  g621(.A(G92gat), .B1(new_n816_), .B2(new_n411_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n469_), .A3(new_n761_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1337gat));
  OAI21_X1  g624(.A(G99gat), .B1(new_n816_), .B2(new_n719_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n264_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n819_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g628(.A1(new_n820_), .A2(new_n499_), .A3(new_n360_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n743_), .A2(new_n360_), .A3(new_n815_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(G106gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n831_), .B2(G106gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  INV_X1    g636(.A(new_n692_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n558_), .A2(new_n683_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n682_), .B(new_n681_), .C1(new_n555_), .C2(new_n557_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n692_), .A2(new_n841_), .A3(KEYINPUT54), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n551_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n654_), .A2(new_n528_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n444_), .B1(new_n846_), .B2(new_n524_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n541_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n846_), .A2(KEYINPUT55), .A3(new_n444_), .A4(new_n524_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n845_), .B1(new_n851_), .B2(new_n545_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n845_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n546_), .B(new_n853_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n844_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n551_), .A2(new_n553_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n588_), .A2(new_n598_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n615_), .B1(new_n607_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n856_), .A2(new_n616_), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n690_), .B1(new_n855_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n524_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n848_), .B1(new_n865_), .B2(new_n445_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n541_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n850_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n545_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n853_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n851_), .A2(new_n545_), .A3(new_n845_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n871_), .A2(new_n617_), .A3(new_n551_), .A4(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n856_), .A2(new_n616_), .A3(new_n860_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n672_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT57), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT121), .B1(new_n877_), .B2(KEYINPUT58), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n551_), .A2(new_n616_), .A3(new_n860_), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT56), .B(new_n546_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n870_), .A2(KEYINPUT56), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n551_), .A2(new_n616_), .A3(new_n860_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n851_), .A2(new_n886_), .A3(new_n545_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n882_), .A4(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n877_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n883_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n736_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n864_), .B(new_n876_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n843_), .B1(new_n893_), .B2(new_n641_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n761_), .A2(new_n360_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n318_), .A3(new_n264_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(G113gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n617_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n889_), .A2(new_n890_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n883_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n892_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n864_), .A2(new_n876_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n641_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n843_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n896_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(KEYINPUT59), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n911_), .A2(new_n683_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n899_), .B1(new_n912_), .B2(new_n898_), .ZN(G1340gat));
  INV_X1    g712(.A(new_n911_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G120gat), .B1(new_n914_), .B2(new_n785_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n897_), .ZN(new_n916_));
  INV_X1    g715(.A(G120gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(KEYINPUT60), .B2(new_n917_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n915_), .B1(new_n916_), .B2(new_n919_), .ZN(G1341gat));
  INV_X1    g719(.A(G127gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n911_), .B2(new_n640_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n916_), .A2(G127gat), .A3(new_n641_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(KEYINPUT123), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1342gat));
  OAI21_X1  g728(.A(G134gat), .B1(new_n914_), .B2(new_n892_), .ZN(new_n930_));
  OR3_X1    g729(.A1(new_n916_), .A2(G134gat), .A3(new_n690_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1343gat));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n264_), .A2(new_n761_), .A3(new_n319_), .A4(new_n361_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n894_), .B2(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n875_), .B(new_n863_), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT58), .B1(new_n888_), .B2(new_n877_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n736_), .B1(new_n938_), .B2(new_n883_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n640_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT124), .B(new_n934_), .C1(new_n940_), .C2(new_n843_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n936_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n617_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n686_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g745(.A(KEYINPUT124), .B1(new_n906_), .B2(new_n934_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n894_), .A2(new_n933_), .A3(new_n935_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n640_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n942_), .A2(KEYINPUT125), .A3(new_n640_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT61), .B(G155gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n953_), .ZN(new_n955_));
  AOI21_X1  g754(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n640_), .ZN(new_n956_));
  AOI211_X1 g755(.A(new_n950_), .B(new_n641_), .C1(new_n936_), .C2(new_n941_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n954_), .A2(new_n958_), .ZN(G1346gat));
  INV_X1    g758(.A(new_n942_), .ZN(new_n960_));
  OR3_X1    g759(.A1(new_n960_), .A2(G162gat), .A3(new_n690_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G162gat), .B1(new_n960_), .B2(new_n892_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n894_), .A2(new_n411_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n719_), .A2(new_n318_), .A3(new_n360_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n966_), .A2(new_n618_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT22), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n969_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n971_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n211_), .B1(new_n967_), .B2(new_n971_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n970_), .B1(new_n972_), .B2(new_n973_), .ZN(G1348gat));
  OAI21_X1  g773(.A(G176gat), .B1(new_n966_), .B2(new_n785_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n558_), .A2(new_n212_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n966_), .B2(new_n976_), .ZN(G1349gat));
  OAI21_X1  g776(.A(new_n223_), .B1(new_n966_), .B2(new_n641_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n370_), .ZN(new_n979_));
  NAND4_X1  g778(.A1(new_n964_), .A2(new_n979_), .A3(new_n640_), .A4(new_n965_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n978_), .B1(KEYINPUT126), .B2(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(KEYINPUT126), .B2(new_n980_), .ZN(G1350gat));
  OAI21_X1  g781(.A(G190gat), .B1(new_n966_), .B2(new_n892_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n672_), .A2(new_n371_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n966_), .B2(new_n984_), .ZN(G1351gat));
  NOR2_X1   g784(.A1(new_n264_), .A2(new_n413_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n964_), .A2(new_n986_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n987_), .A2(new_n618_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(new_n336_), .ZN(G1352gat));
  NOR2_X1   g788(.A1(new_n987_), .A2(new_n785_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(new_n333_), .ZN(G1353gat));
  INV_X1    g790(.A(new_n987_), .ZN(new_n992_));
  XOR2_X1   g791(.A(KEYINPUT63), .B(G211gat), .Z(new_n993_));
  NAND3_X1  g792(.A1(new_n992_), .A2(new_n640_), .A3(new_n993_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n994_), .A2(KEYINPUT127), .ZN(new_n995_));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996_));
  NAND4_X1  g795(.A1(new_n992_), .A2(new_n996_), .A3(new_n640_), .A4(new_n993_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n998_), .B1(new_n987_), .B2(new_n641_), .ZN(new_n999_));
  AND3_X1   g798(.A1(new_n995_), .A2(new_n997_), .A3(new_n999_), .ZN(G1354gat));
  OAI21_X1  g799(.A(G218gat), .B1(new_n987_), .B2(new_n892_), .ZN(new_n1001_));
  OR2_X1    g800(.A1(new_n690_), .A2(G218gat), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n987_), .B2(new_n1002_), .ZN(G1355gat));
endmodule


