//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n206_), .A2(new_n207_), .A3(new_n204_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n215_), .A3(KEYINPUT86), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT77), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n232_), .B2(new_n228_), .ZN(new_n233_));
  AND2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT78), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT23), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT79), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n235_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n233_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n244_), .A3(KEYINPUT23), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  INV_X1    g050(.A(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n231_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT22), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(G169gat), .ZN(new_n257_));
  INV_X1    g056(.A(G169gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT22), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G176gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n255_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n227_), .A2(new_n247_), .B1(new_n254_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n203_), .B1(new_n220_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT23), .B1(new_n242_), .B2(new_n244_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n253_), .B1(new_n265_), .B2(new_n239_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT89), .B1(new_n257_), .B2(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n258_), .A2(KEYINPUT22), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(G169gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT89), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n261_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n266_), .A2(new_n272_), .A3(new_n231_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(G183gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n251_), .A2(KEYINPUT25), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT88), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n251_), .A2(KEYINPUT25), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(G183gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n222_), .A3(new_n281_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n232_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n228_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n250_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n273_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n216_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n264_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n212_), .A2(new_n215_), .A3(KEYINPUT86), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT86), .B1(new_n212_), .B2(new_n215_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT77), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT77), .B1(new_n221_), .B2(new_n222_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n286_), .B1(new_n265_), .B2(new_n239_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n248_), .A2(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n260_), .A2(new_n261_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n231_), .ZN(new_n303_));
  OAI22_X1  g102(.A1(new_n299_), .A2(new_n300_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n292_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n212_), .A2(new_n215_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n273_), .A2(new_n287_), .A3(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n305_), .A2(KEYINPUT20), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n293_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n293_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT27), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n319_), .A3(KEYINPUT20), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n305_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n308_), .B2(KEYINPUT20), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n292_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n220_), .A2(new_n263_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n324_), .A2(new_n289_), .A3(KEYINPUT20), .A4(new_n306_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT96), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n264_), .A2(KEYINPUT96), .A3(new_n306_), .A4(new_n289_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n314_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT99), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(KEYINPUT99), .A3(new_n314_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n317_), .A2(KEYINPUT27), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n318_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n351_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT82), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G155gat), .ZN(new_n361_));
  INV_X1    g160(.A(G162gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n345_), .B1(new_n357_), .B2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n360_), .A2(new_n366_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n352_), .A2(new_n353_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT2), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n350_), .A4(new_n349_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n373_), .A3(KEYINPUT83), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n352_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n365_), .A2(KEYINPUT1), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n359_), .B1(new_n358_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n344_), .B1(new_n375_), .B2(new_n383_), .ZN(new_n384_));
  AOI211_X1 g183(.A(new_n343_), .B(new_n382_), .C1(new_n368_), .C2(new_n374_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT4), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n343_), .A2(KEYINPUT4), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n369_), .A2(KEYINPUT83), .A3(new_n373_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT83), .B1(new_n369_), .B2(new_n373_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n383_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n386_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n397_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT92), .B(new_n397_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n399_), .A2(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n386_), .A2(new_n396_), .A3(KEYINPUT91), .A4(new_n398_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n340_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT90), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n394_), .B1(new_n393_), .B2(new_n388_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n393_), .A2(new_n343_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n387_), .A2(new_n344_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n400_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n403_), .A2(new_n404_), .ZN(new_n416_));
  AND4_X1   g215(.A1(new_n340_), .A2(new_n415_), .A3(new_n406_), .A4(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n407_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n383_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G22gat), .B(G50gat), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n387_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n420_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n426_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT85), .A3(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G228gat), .A2(G233gat), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n437_), .B(new_n296_), .C1(new_n387_), .C2(new_n421_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n307_), .B1(new_n393_), .B2(KEYINPUT29), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n437_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n438_), .B(new_n441_), .C1(new_n439_), .C2(new_n437_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n419_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n430_), .A2(new_n435_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT87), .A3(new_n444_), .A4(new_n443_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n434_), .A3(new_n433_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n336_), .A2(new_n418_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n293_), .A2(new_n309_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n314_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT94), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n329_), .A2(KEYINPUT97), .A3(new_n455_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT97), .B1(new_n329_), .B2(new_n455_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(new_n418_), .B2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n453_), .A2(new_n456_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n329_), .A2(new_n455_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n466_), .B2(new_n458_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n415_), .A2(new_n406_), .A3(new_n416_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n340_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n405_), .A2(new_n340_), .A3(new_n406_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n472_), .A3(KEYINPUT98), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n386_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT93), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n398_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n469_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n315_), .A2(new_n479_), .A3(new_n317_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n471_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n462_), .A2(new_n473_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n450_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n451_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n263_), .B(KEYINPUT30), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(G15gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G71gat), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n488_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n343_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT80), .B(G43gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT31), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n496_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n202_), .B1(new_n487_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n467_), .A2(new_n472_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n502_), .A2(new_n452_), .B1(new_n483_), .B2(new_n482_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n450_), .B1(new_n503_), .B2(new_n473_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT100), .B(new_n499_), .C1(new_n504_), .C2(new_n451_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n336_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(new_n450_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n507_), .A3(new_n418_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G43gat), .B(G50gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT15), .Z(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT74), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(KEYINPUT74), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n513_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n512_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n522_), .B(new_n512_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G113gat), .B(G141gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n530_), .B(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n509_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT6), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT65), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(KEYINPUT65), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(KEYINPUT6), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(G99gat), .A4(G106gat), .ZN(new_n544_));
  INV_X1    g343(.A(G106gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n493_), .A2(new_n545_), .A3(KEYINPUT66), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT7), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(new_n493_), .A3(new_n545_), .A4(KEYINPUT66), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n541_), .A2(new_n544_), .A3(new_n547_), .A4(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT8), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G85gat), .B(G92gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(KEYINPUT67), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n541_), .A2(new_n544_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT10), .B(G99gat), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n545_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT64), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(KEYINPUT64), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n551_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n560_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n557_), .A2(new_n559_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n555_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n568_), .A2(new_n512_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n572_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT72), .Z(new_n575_));
  NOR2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n565_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n550_), .A2(new_n551_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n555_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT69), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n556_), .A2(new_n582_), .A3(new_n567_), .A4(new_n565_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n513_), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n576_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT71), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n573_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n574_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT73), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT36), .Z(new_n596_));
  INV_X1    g395(.A(KEYINPUT73), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n574_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n585_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G120gat), .B(G148gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n563_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n541_), .A2(new_n544_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n580_), .A2(new_n612_), .A3(new_n566_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G71gat), .B(G78gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G57gat), .B(G64gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(KEYINPUT11), .B2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(KEYINPUT11), .B2(new_n615_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n614_), .A3(KEYINPUT11), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n568_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n609_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT68), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(KEYINPUT12), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n581_), .A2(new_n583_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT12), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n613_), .B2(new_n619_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n628_), .A2(new_n609_), .A3(new_n620_), .A4(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n608_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n631_), .A3(new_n608_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(KEYINPUT13), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT13), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n623_), .A2(KEYINPUT68), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n623_), .A2(KEYINPUT68), .ZN(new_n638_));
  AND4_X1   g437(.A1(new_n631_), .A2(new_n637_), .A3(new_n638_), .A4(new_n608_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n632_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n596_), .B1(new_n598_), .B2(new_n585_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n602_), .A2(KEYINPUT37), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT17), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n648_), .A2(KEYINPUT75), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n522_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n621_), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n650_), .B(new_n653_), .C1(new_n649_), .C2(new_n648_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(new_n650_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n603_), .A2(new_n641_), .A3(new_n643_), .A4(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n535_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n514_), .A3(new_n472_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT101), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n661_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT102), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n600_), .A2(new_n602_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n509_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n641_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n534_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n657_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G1gat), .B1(new_n671_), .B2(new_n418_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n663_), .A2(new_n665_), .A3(new_n672_), .ZN(G1324gat));
  NAND3_X1  g472(.A1(new_n659_), .A2(new_n515_), .A3(new_n506_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n506_), .A3(new_n670_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n515_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT40), .B(new_n674_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1325gat));
  NAND3_X1  g485(.A1(new_n659_), .A2(new_n490_), .A3(new_n500_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n667_), .A2(new_n500_), .A3(new_n670_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT104), .Z(G1326gat));
  OAI21_X1  g491(.A(G22gat), .B1(new_n671_), .B2(new_n486_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n486_), .A2(G22gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT106), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n659_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n509_), .A2(new_n534_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n666_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n657_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n700_), .A2(new_n641_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G29gat), .B1(new_n703_), .B2(new_n472_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n669_), .A2(new_n656_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT37), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n643_), .B1(new_n666_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n509_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT43), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n509_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n706_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT107), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n715_));
  INV_X1    g514(.A(new_n713_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n509_), .B2(new_n709_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n705_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n705_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n723_), .A2(G29gat), .A3(new_n472_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n704_), .B1(new_n722_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n506_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n722_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n703_), .A2(new_n727_), .A3(new_n506_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT45), .Z(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n731_), .B(KEYINPUT45), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n728_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT46), .B(new_n734_), .C1(new_n735_), .C2(new_n727_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1329gat));
  AND2_X1   g536(.A1(new_n703_), .A2(new_n500_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(G43gat), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n715_), .A2(new_n721_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n723_), .A2(G43gat), .A3(new_n500_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n740_), .B(new_n741_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n741_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n739_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1330gat));
  AOI21_X1  g547(.A(G50gat), .B1(new_n703_), .B2(new_n450_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n723_), .A2(G50gat), .A3(new_n450_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n722_), .B2(new_n750_), .ZN(G1331gat));
  INV_X1    g550(.A(new_n534_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n667_), .A2(new_n752_), .A3(new_n656_), .A4(new_n641_), .ZN(new_n753_));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n418_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n509_), .A2(new_n752_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n709_), .A2(new_n657_), .A3(new_n668_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n418_), .B1(new_n759_), .B2(KEYINPUT109), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(KEYINPUT109), .B2(new_n759_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n761_), .B2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g561(.A(G64gat), .B1(new_n753_), .B2(new_n336_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT48), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n336_), .A2(G64gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n758_), .B2(new_n765_), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n753_), .B2(new_n499_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT49), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n499_), .A2(G71gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n758_), .B2(new_n769_), .ZN(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n753_), .B2(new_n486_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT50), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n486_), .A2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n758_), .B2(new_n773_), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n702_), .A2(new_n668_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n756_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(G85gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n472_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n668_), .A2(new_n534_), .A3(new_n656_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT110), .Z(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n472_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n782_), .B2(new_n777_), .ZN(G1336gat));
  AOI21_X1  g582(.A(G92gat), .B1(new_n776_), .B2(new_n506_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n506_), .A2(G92gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT111), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n781_), .B2(new_n786_), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n776_), .A2(new_n500_), .A3(new_n558_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT112), .ZN(new_n789_));
  OAI21_X1  g588(.A(G99gat), .B1(new_n780_), .B2(new_n499_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT51), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n776_), .A2(new_n545_), .A3(new_n450_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n450_), .B(new_n779_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g601(.A(new_n526_), .B1(new_n525_), .B2(KEYINPUT117), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(KEYINPUT117), .B2(new_n525_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n533_), .B1(new_n529_), .B2(new_n526_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n530_), .A2(new_n533_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n634_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n631_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n609_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n628_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n630_), .A2(new_n620_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n577_), .A2(new_n580_), .A3(new_n621_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n622_), .B2(new_n629_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n815_), .A2(KEYINPUT55), .A3(new_n609_), .A4(new_n628_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(new_n813_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT115), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n809_), .A2(new_n813_), .A3(new_n816_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n607_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n823_), .B(new_n608_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n807_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT58), .B(new_n807_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n827_), .A2(new_n709_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n821_), .A2(new_n607_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n823_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n607_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n534_), .A2(new_n634_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n824_), .B2(KEYINPUT116), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n633_), .A2(new_n634_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n834_), .A2(new_n836_), .B1(new_n837_), .B2(new_n806_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n701_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n806_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n822_), .A2(new_n824_), .A3(KEYINPUT116), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n534_), .B(new_n634_), .C1(new_n833_), .C2(new_n832_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n666_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n829_), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n656_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n829_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n701_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n844_), .B1(new_n843_), .B2(new_n666_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n657_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n708_), .A2(new_n668_), .A3(new_n752_), .A4(new_n656_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n854_), .B2(KEYINPUT113), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n658_), .A2(new_n856_), .A3(new_n857_), .A4(new_n752_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(KEYINPUT113), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n855_), .A2(new_n858_), .A3(new_n861_), .A4(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n847_), .A2(new_n853_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n500_), .A2(new_n507_), .A3(new_n472_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n752_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n851_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n846_), .A2(KEYINPUT118), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n657_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n868_), .B1(new_n876_), .B2(new_n865_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n870_), .B(new_n872_), .C1(new_n877_), .C2(new_n867_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n875_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n657_), .B1(new_n846_), .B2(KEYINPUT118), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n865_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n534_), .A3(new_n869_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n871_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n878_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n878_), .A2(KEYINPUT120), .A3(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1340gat));
  XOR2_X1   g687(.A(KEYINPUT121), .B(G120gat), .Z(new_n889_));
  OR2_X1    g688(.A1(new_n889_), .A2(KEYINPUT60), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n668_), .B2(KEYINPUT60), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n881_), .A2(new_n869_), .A3(new_n890_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n870_), .B1(new_n877_), .B2(new_n867_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n668_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n889_), .B2(new_n896_), .ZN(G1341gat));
  OAI21_X1  g696(.A(G127gat), .B1(new_n895_), .B2(new_n657_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n877_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n657_), .A2(G127gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n895_), .B2(new_n708_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n666_), .A2(G134gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n899_), .B2(new_n903_), .ZN(G1343gat));
  AOI21_X1  g703(.A(new_n500_), .B1(new_n876_), .B2(new_n865_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n506_), .A2(new_n486_), .A3(new_n418_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n752_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT123), .B(G141gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n668_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n348_), .ZN(G1345gat));
  NOR2_X1   g711(.A1(new_n907_), .A2(new_n657_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT61), .B(G155gat), .Z(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n907_), .B2(new_n708_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n701_), .A2(new_n362_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n907_), .B2(new_n917_), .ZN(G1347gat));
  NOR4_X1   g717(.A1(new_n499_), .A2(new_n472_), .A3(new_n450_), .A4(new_n336_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n866_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n534_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(G169gat), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n920_), .A2(new_n534_), .A3(new_n267_), .A4(new_n271_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1348gat));
  AND2_X1   g726(.A1(new_n881_), .A2(new_n919_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n668_), .A2(new_n261_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n928_), .A2(KEYINPUT124), .A3(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT124), .B1(new_n928_), .B2(new_n929_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G176gat), .B1(new_n920_), .B2(new_n641_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(G1349gat));
  NAND2_X1  g732(.A1(new_n866_), .A2(new_n919_), .ZN(new_n934_));
  AOI211_X1 g733(.A(new_n657_), .B(new_n934_), .C1(new_n277_), .C2(new_n281_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n928_), .A2(new_n656_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937_));
  AOI21_X1  g736(.A(G183gat), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n928_), .A2(KEYINPUT125), .A3(new_n656_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n920_), .A2(new_n222_), .A3(new_n701_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G190gat), .B1(new_n934_), .B2(new_n708_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(new_n942_), .A3(KEYINPUT126), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n486_), .A2(new_n336_), .A3(new_n472_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n905_), .A2(new_n534_), .A3(new_n948_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g749(.A1(new_n905_), .A2(new_n641_), .A3(new_n948_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g751(.A(new_n657_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n905_), .A2(new_n948_), .A3(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT127), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n954_), .B(new_n956_), .ZN(G1354gat));
  NAND2_X1  g756(.A1(new_n905_), .A2(new_n948_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G218gat), .B1(new_n958_), .B2(new_n708_), .ZN(new_n959_));
  INV_X1    g758(.A(G218gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n701_), .A2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n959_), .B1(new_n958_), .B2(new_n961_), .ZN(G1355gat));
endmodule


