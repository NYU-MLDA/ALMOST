//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  AND2_X1   g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT72), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT70), .B(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT71), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G1gat), .B(G8gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n216_), .B(KEYINPUT71), .ZN(new_n221_));
  INV_X1    g020(.A(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n211_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT74), .ZN(new_n227_));
  XOR2_X1   g026(.A(G127gat), .B(G155gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT17), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n227_), .B(new_n233_), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n226_), .A2(KEYINPUT17), .A3(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT75), .Z(new_n237_));
  XOR2_X1   g036(.A(G85gat), .B(G92gat), .Z(new_n238_));
  NOR2_X1   g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT7), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G99gat), .A2(G106gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT6), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n238_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT8), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT64), .B(G106gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT65), .ZN(new_n250_));
  INV_X1    g049(.A(G85gat), .ZN(new_n251_));
  INV_X1    g050(.A(G92gat), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n251_), .A2(new_n252_), .A3(KEYINPUT9), .ZN(new_n253_));
  AOI211_X1 g052(.A(new_n253_), .B(new_n244_), .C1(KEYINPUT9), .C2(new_n238_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n246_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G29gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT15), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n246_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G232gat), .A2(G233gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT34), .Z(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT66), .B(KEYINPUT35), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI211_X1 g068(.A(new_n266_), .B(new_n265_), .C1(new_n261_), .C2(KEYINPUT67), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n263_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G134gat), .B(G162gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT69), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT37), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n256_), .B(new_n208_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT12), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n208_), .B1(new_n246_), .B2(new_n255_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G230gat), .A2(G233gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n287_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G120gat), .B(G148gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT5), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G176gat), .B(G204gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n295_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT13), .Z(new_n305_));
  NOR3_X1   g104(.A1(new_n237_), .A2(new_n286_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n224_), .A2(new_n259_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT76), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n307_), .B2(KEYINPUT76), .ZN(new_n311_));
  OAI22_X1  g110(.A1(new_n310_), .A2(new_n311_), .B1(new_n259_), .B2(new_n224_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n224_), .A2(new_n259_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n225_), .A2(new_n260_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n316_), .A3(new_n307_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G169gat), .B(G197gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n330_), .ZN(new_n333_));
  INV_X1    g132(.A(G169gat), .ZN(new_n334_));
  INV_X1    g133(.A(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT24), .A3(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n333_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G183gat), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT78), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G190gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n347_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n330_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n332_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n352_), .A3(new_n344_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G169gat), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n343_), .A2(new_n355_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G71gat), .B(G99gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(G15gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n367_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(G134gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G127gat), .ZN(new_n374_));
  INV_X1    g173(.A(G127gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G120gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G113gat), .ZN(new_n379_));
  INV_X1    g178(.A(G113gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G120gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n377_), .B2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n374_), .A2(new_n376_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n379_), .A2(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n388_), .B2(KEYINPUT80), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT31), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n372_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394_));
  OR3_X1    g193(.A1(new_n372_), .A2(new_n394_), .A3(new_n390_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n372_), .B2(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT19), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n358_), .B1(new_n332_), .B2(new_n356_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n348_), .A2(new_n349_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n345_), .B(new_n346_), .C1(new_n402_), .C2(new_n354_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT24), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n340_), .A2(KEYINPUT92), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n336_), .B(new_n337_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n339_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n401_), .A2(new_n403_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n363_), .B1(new_n333_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G218gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G211gat), .ZN(new_n415_));
  INV_X1    g214(.A(G211gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G218gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G197gat), .A2(G204gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G197gat), .A2(G204gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT21), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT21), .ZN(new_n422_));
  AND2_X1   g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G197gat), .A2(G204gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n422_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT89), .B1(new_n423_), .B2(new_n424_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n430_), .A3(new_n420_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT90), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT90), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n428_), .A2(new_n431_), .A3(new_n429_), .A4(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n427_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n364_), .A2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n400_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G8gat), .B(G36gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT18), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n433_), .A2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n426_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n343_), .A2(new_n355_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n361_), .A2(new_n363_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n400_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n426_), .A3(new_n412_), .A4(new_n410_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(KEYINPUT20), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n439_), .A2(new_n443_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n443_), .B1(new_n439_), .B2(new_n452_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n456_));
  OR3_X1    g255(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462_));
  INV_X1    g261(.A(G155gat), .ZN(new_n463_));
  INV_X1    g262(.A(G162gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n465_), .A2(new_n466_), .B1(KEYINPUT1), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT1), .ZN(new_n469_));
  INV_X1    g268(.A(new_n467_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n468_), .A2(KEYINPUT85), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(KEYINPUT1), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n461_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G141gat), .A2(G148gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT3), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n460_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n481_), .A2(new_n483_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n470_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n388_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n456_), .B1(new_n477_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n389_), .B1(new_n477_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n461_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n472_), .A2(KEYINPUT85), .A3(new_n473_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n470_), .A2(new_n469_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n468_), .A2(KEYINPUT85), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n487_), .A2(new_n488_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(KEYINPUT93), .A3(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT4), .A4(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n377_), .A2(new_n382_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n374_), .A2(new_n376_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT80), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n383_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n499_), .B2(new_n489_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n504_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n502_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n502_), .A2(new_n512_), .A3(KEYINPUT94), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G29gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n251_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT0), .B(G57gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n491_), .A2(new_n493_), .A3(new_n501_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n504_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n502_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n491_), .A2(new_n493_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n520_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n502_), .A2(new_n525_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n520_), .A2(KEYINPUT33), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n455_), .A2(new_n523_), .A3(new_n529_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT95), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n439_), .A2(new_n452_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n443_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n439_), .A2(new_n443_), .A3(new_n452_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n537_), .A2(new_n532_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n523_), .A4(new_n529_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n530_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n520_), .B1(new_n530_), .B2(new_n527_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(KEYINPUT98), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n545_), .B(new_n520_), .C1(new_n530_), .C2(new_n527_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n439_), .A2(new_n452_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n410_), .A2(new_n412_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n445_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n364_), .A2(new_n436_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n551_), .A2(KEYINPUT20), .A3(new_n552_), .A4(new_n450_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n451_), .B(KEYINPUT20), .C1(new_n364_), .C2(new_n436_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n553_), .A2(KEYINPUT96), .B1(new_n554_), .B2(new_n400_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n445_), .B2(new_n550_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n450_), .A4(new_n552_), .ZN(new_n559_));
  AOI211_X1 g358(.A(KEYINPUT97), .B(new_n548_), .C1(new_n555_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(KEYINPUT96), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n400_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n548_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n549_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n534_), .B(new_n541_), .C1(new_n547_), .C2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT91), .B(G106gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n571_));
  INV_X1    g370(.A(G228gat), .ZN(new_n572_));
  INV_X1    g371(.A(G233gat), .ZN(new_n573_));
  OAI22_X1  g372(.A1(new_n436_), .A2(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G22gat), .B(G50gat), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  OAI221_X1 g376(.A(new_n577_), .B1(new_n572_), .B2(new_n573_), .C1(new_n436_), .C2(new_n571_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n499_), .A2(new_n489_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(KEYINPUT29), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n477_), .A2(new_n492_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n584_));
  INV_X1    g383(.A(new_n580_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n579_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n576_), .A2(new_n582_), .A3(new_n578_), .A4(new_n586_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n584_), .B1(new_n499_), .B2(new_n489_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G78gat), .B1(new_n590_), .B2(new_n436_), .ZN(new_n591_));
  INV_X1    g390(.A(G78gat), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n445_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n570_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n569_), .A3(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT27), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n453_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n564_), .A2(new_n536_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n537_), .A2(new_n538_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n604_), .A2(new_n605_), .B1(new_n606_), .B2(new_n603_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(new_n547_), .A3(new_n598_), .A4(new_n600_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n568_), .A2(new_n601_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n598_), .A2(new_n600_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n610_), .A2(KEYINPUT99), .A3(new_n547_), .A4(new_n607_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n398_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  INV_X1    g412(.A(new_n607_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n398_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n547_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n612_), .A2(new_n613_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n534_), .A2(new_n541_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n567_), .A2(new_n547_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n601_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n608_), .A2(new_n602_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n611_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT100), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n329_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n306_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n212_), .B1(KEYINPUT101), .B2(KEYINPUT38), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n628_), .A2(new_n547_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT101), .A2(KEYINPUT38), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n618_), .A2(new_n615_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n284_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n305_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(KEYINPUT102), .A3(new_n328_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n305_), .B2(new_n329_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n236_), .A3(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n639_), .A2(new_n547_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G1gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n632_), .B1(new_n645_), .B2(new_n646_), .ZN(G1324gat));
  NAND4_X1  g446(.A1(new_n306_), .A2(new_n627_), .A3(new_n213_), .A4(new_n614_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n644_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(new_n614_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G8gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G8gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  NOR2_X1   g455(.A1(new_n639_), .A2(new_n644_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n369_), .B1(new_n657_), .B2(new_n398_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n628_), .A2(G15gat), .A3(new_n616_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT104), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(G1326gat));
  OR3_X1    g463(.A1(new_n628_), .A2(G22gat), .A3(new_n601_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n657_), .A2(new_n610_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  XNOR2_X1  g469(.A(new_n236_), .B(KEYINPUT75), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n284_), .A3(new_n305_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n627_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G29gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n617_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n641_), .A2(new_n237_), .A3(new_n643_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT43), .B(new_n285_), .C1(new_n619_), .C2(new_n626_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n635_), .B2(new_n286_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n678_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n634_), .A2(new_n633_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n612_), .A2(new_n613_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n286_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n635_), .A2(new_n680_), .A3(new_n286_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n689_), .B2(new_n678_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n683_), .A2(new_n690_), .A3(new_n547_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n676_), .B1(new_n691_), .B2(new_n675_), .ZN(G1328gat));
  OR2_X1    g491(.A1(new_n614_), .A2(KEYINPUT106), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n614_), .A2(KEYINPUT106), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n673_), .A2(G36gat), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n678_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n614_), .A3(new_n682_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(KEYINPUT105), .A3(new_n614_), .A4(new_n682_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT46), .B(new_n699_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n706_), .A2(G36gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n704_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n698_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1329gat));
  AOI21_X1  g512(.A(G43gat), .B1(new_n674_), .B2(new_n398_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n683_), .A2(new_n690_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n398_), .A2(G43gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1330gat));
  OR3_X1    g518(.A1(new_n673_), .A2(G50gat), .A3(new_n601_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n715_), .A2(new_n610_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT109), .B1(new_n721_), .B2(G50gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  NOR2_X1   g523(.A1(new_n640_), .A2(new_n328_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n635_), .A2(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(new_n671_), .A3(new_n285_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n617_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n725_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n639_), .A2(new_n237_), .A3(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n617_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n732_), .B2(new_n728_), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n727_), .A2(new_n734_), .A3(new_n695_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(new_n695_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G64gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT48), .B(new_n734_), .C1(new_n731_), .C2(new_n695_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n398_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT110), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n727_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n731_), .A2(new_n398_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G71gat), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT49), .B(new_n741_), .C1(new_n731_), .C2(new_n398_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  NAND3_X1  g548(.A1(new_n727_), .A2(new_n592_), .A3(new_n610_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n731_), .A2(new_n610_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G78gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT50), .B(new_n592_), .C1(new_n731_), .C2(new_n610_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(G1335gat));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n689_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n730_), .A2(new_n671_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n687_), .A2(KEYINPUT111), .A3(new_n688_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n547_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n284_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n726_), .A2(new_n762_), .A3(new_n237_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n251_), .A3(new_n617_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n696_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n252_), .A3(new_n614_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n760_), .B2(new_n616_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(new_n247_), .A3(new_n398_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n763_), .A2(new_n248_), .A3(new_n610_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n689_), .A2(new_n610_), .A3(new_n758_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND4_X1   g575(.A1(KEYINPUT113), .A2(new_n775_), .A3(new_n776_), .A4(G106gat), .ZN(new_n777_));
  INV_X1    g576(.A(G106gat), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(KEYINPUT52), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n775_), .A2(new_n780_), .B1(KEYINPUT113), .B2(new_n776_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n774_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n616_), .A2(new_n547_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n615_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n316_), .B1(new_n224_), .B2(new_n259_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n324_), .B1(new_n319_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n327_), .A2(new_n303_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n293_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n288_), .A2(new_n791_), .A3(new_n291_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(KEYINPUT55), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n294_), .B2(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n793_), .A2(KEYINPUT116), .A3(new_n796_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n794_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n300_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n790_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n292_), .A2(KEYINPUT55), .A3(new_n293_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n288_), .A2(new_n791_), .A3(new_n291_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT116), .B1(new_n793_), .B2(new_n796_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n294_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n810_), .B2(new_n302_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n300_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT118), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n803_), .A2(new_n813_), .A3(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT119), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n803_), .A2(new_n813_), .A3(new_n816_), .A4(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT58), .B1(new_n803_), .B2(new_n813_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n285_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n823_), .A3(new_n820_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n810_), .B2(new_n302_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n804_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(KEYINPUT56), .C1(new_n810_), .C2(new_n302_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n328_), .A3(new_n303_), .A4(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n304_), .A2(new_n327_), .A3(new_n789_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n831_), .B2(new_n284_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n762_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(new_n824_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n236_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT114), .B1(new_n237_), .B2(new_n328_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n671_), .A2(new_n840_), .A3(new_n329_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n286_), .A2(new_n305_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT54), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n785_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n328_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(new_n844_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n785_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n671_), .B1(new_n835_), .B2(new_n821_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n844_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n848_), .A2(new_n853_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n849_), .A2(KEYINPUT59), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n380_), .B1(new_n328_), .B2(KEYINPUT122), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(KEYINPUT122), .B2(new_n380_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n846_), .B1(new_n855_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n843_), .B(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n854_), .B1(new_n860_), .B2(new_n850_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n305_), .B(new_n861_), .C1(new_n845_), .C2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n378_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n378_), .A2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(KEYINPUT123), .B2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n845_), .B(new_n867_), .C1(KEYINPUT123), .C2(new_n865_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n845_), .B2(new_n671_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n236_), .A2(G127gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT124), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n855_), .B2(new_n872_), .ZN(G1342gat));
  OAI211_X1 g672(.A(new_n286_), .B(new_n861_), .C1(new_n845_), .C2(new_n862_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G134gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n845_), .A2(new_n373_), .A3(new_n762_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1343gat));
  NOR4_X1   g676(.A1(new_n695_), .A2(new_n547_), .A3(new_n398_), .A4(new_n601_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n847_), .A2(new_n328_), .A3(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g679(.A1(new_n847_), .A2(new_n305_), .A3(new_n878_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g681(.A1(new_n847_), .A2(new_n671_), .A3(new_n878_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  NAND4_X1  g684(.A1(new_n847_), .A2(new_n464_), .A3(new_n762_), .A4(new_n878_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n847_), .A2(new_n286_), .A3(new_n878_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n464_), .ZN(G1347gat));
  XNOR2_X1  g687(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n618_), .A2(new_n695_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n610_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n328_), .B(new_n891_), .C1(new_n860_), .C2(new_n850_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n889_), .B1(new_n892_), .B2(KEYINPUT22), .ZN(new_n893_));
  OAI21_X1  g692(.A(G169gat), .B1(new_n892_), .B2(new_n889_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n334_), .B2(new_n893_), .ZN(G1348gat));
  OAI211_X1 g695(.A(new_n305_), .B(new_n891_), .C1(new_n860_), .C2(new_n850_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT126), .B1(new_n898_), .B2(G176gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n900_), .A3(new_n335_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n610_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n640_), .A2(new_n890_), .A3(new_n335_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n899_), .A2(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NAND4_X1  g703(.A1(new_n902_), .A2(new_n618_), .A3(new_n671_), .A4(new_n695_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n852_), .A2(new_n891_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n837_), .A2(new_n347_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n905_), .A2(new_n344_), .B1(new_n906_), .B2(new_n907_), .ZN(G1350gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n286_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G190gat), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n906_), .B(new_n762_), .C1(new_n354_), .C2(new_n402_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NOR4_X1   g711(.A1(new_n696_), .A2(new_n617_), .A3(new_n398_), .A4(new_n601_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n328_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n305_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n236_), .B1(new_n920_), .B2(new_n416_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n915_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n416_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(new_n915_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G218gat), .B1(new_n926_), .B2(new_n285_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n915_), .A2(new_n414_), .A3(new_n762_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1355gat));
endmodule


