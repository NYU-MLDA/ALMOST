//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  OR2_X1    g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT87), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n202_), .B(new_n203_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n203_), .B(KEYINPUT2), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n202_), .B2(KEYINPUT89), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n202_), .A2(KEYINPUT89), .A3(KEYINPUT3), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n208_), .B(new_n211_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT90), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT28), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n228_), .A3(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G22gat), .B(G50gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n233_));
  AOI211_X1 g032(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n221_), .C2(new_n223_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT21), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n240_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT21), .B1(new_n242_), .B2(new_n243_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n220_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(new_n225_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G228gat), .A3(G233gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n247_), .A2(new_n248_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(G228gat), .B2(G233gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n256_), .A2(KEYINPUT93), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n231_), .A2(new_n235_), .A3(KEYINPUT91), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(KEYINPUT93), .A3(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n238_), .A2(new_n258_), .A3(new_n259_), .A4(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n260_), .A2(new_n231_), .A3(new_n262_), .A4(new_n235_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G183gat), .A3(G190gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT84), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT23), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n275_), .B2(KEYINPUT84), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT83), .B(G176gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT22), .B(G169gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  INV_X1    g084(.A(G183gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT82), .B1(new_n286_), .B2(KEYINPUT25), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT25), .B(G183gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n287_), .C1(new_n288_), .C2(KEYINPUT82), .ZN(new_n289_));
  NOR3_X1   g088(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n292_), .B2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n274_), .A2(new_n271_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n279_), .A2(new_n284_), .B1(new_n289_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n269_), .B1(new_n253_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n283_), .B(KEYINPUT96), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n282_), .B(new_n298_), .C1(new_n275_), .C2(new_n277_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT95), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT94), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n285_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n285_), .A2(new_n302_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n303_), .A2(new_n288_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n276_), .A2(new_n293_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n285_), .B(KEYINPUT94), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n288_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(KEYINPUT95), .A3(new_n293_), .A4(new_n276_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n300_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n297_), .B1(new_n311_), .B2(new_n253_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT19), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n253_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n314_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n296_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n269_), .B1(new_n318_), .B2(new_n249_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G8gat), .B(G36gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n315_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n268_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n297_), .B(new_n317_), .C1(new_n311_), .C2(new_n253_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n299_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT101), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT101), .B(new_n299_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n253_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n317_), .B1(new_n336_), .B2(new_n319_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n325_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n315_), .A2(new_n320_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(KEYINPUT27), .C1(new_n325_), .C2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT103), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n329_), .A2(new_n340_), .A3(KEYINPUT103), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n266_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT86), .Z(new_n349_));
  NAND3_X1  g148(.A1(new_n221_), .A2(new_n349_), .A3(new_n223_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n250_), .A2(new_n348_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT4), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n221_), .A2(new_n349_), .A3(new_n355_), .A4(new_n223_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G1gat), .B(G29gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n358_), .A2(new_n364_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n359_), .A2(new_n365_), .B1(new_n366_), .B2(new_n357_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n296_), .B(KEYINPUT30), .Z(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT85), .B(G43gat), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(G15gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G71gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n349_), .B(KEYINPUT31), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G99gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n373_), .A2(new_n376_), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n368_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n345_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n329_), .A2(new_n367_), .A3(new_n340_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n265_), .B2(new_n264_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n366_), .A2(new_n357_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT99), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(KEYINPUT99), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n327_), .A2(new_n328_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT100), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n352_), .A2(KEYINPUT100), .A3(new_n353_), .A4(new_n356_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n350_), .A2(new_n351_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n364_), .B1(new_n400_), .B2(new_n354_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n339_), .B2(new_n404_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n394_), .A2(new_n403_), .B1(new_n367_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n266_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n388_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n383_), .A2(new_n384_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n386_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G190gat), .B(G218gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT77), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G134gat), .B(G162gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT36), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT15), .ZN(new_n417_));
  INV_X1    g216(.A(G50gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G43gat), .ZN(new_n419_));
  INV_X1    g218(.A(G43gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G50gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G29gat), .B(G36gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G36gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G29gat), .ZN(new_n426_));
  INV_X1    g225(.A(G29gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G36gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n424_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n424_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n417_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n432_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n429_), .A2(new_n430_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n422_), .A2(new_n423_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n424_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT15), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT65), .B(G106gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT64), .B1(new_n452_), .B2(new_n445_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n444_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n455_), .A2(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G85gat), .ZN(new_n460_));
  INV_X1    g259(.A(G92gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT67), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n462_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n454_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT68), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n448_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n452_), .A2(KEYINPUT64), .A3(new_n445_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n479_), .B2(new_n444_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n467_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n474_), .A2(new_n475_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n474_), .B2(new_n482_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n472_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT69), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n451_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G85gat), .B(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n487_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n494_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n487_), .B(new_n498_), .C1(new_n476_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n486_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT69), .B1(new_n469_), .B2(new_n471_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n497_), .B1(new_n505_), .B2(new_n490_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT70), .B(new_n501_), .C1(new_n506_), .C2(new_n487_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n443_), .B1(new_n485_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n501_), .B1(new_n506_), .B2(new_n487_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(new_n482_), .A3(new_n474_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n439_), .A2(new_n440_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n509_), .A2(KEYINPUT76), .A3(new_n515_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n473_), .A2(KEYINPUT68), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n481_), .B1(new_n480_), .B2(new_n467_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT71), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n474_), .A2(new_n475_), .A3(new_n482_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n503_), .A2(new_n507_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n442_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n520_), .B1(new_n527_), .B2(new_n514_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n526_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n514_), .B1(new_n530_), .B2(new_n443_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n518_), .B1(new_n531_), .B2(KEYINPUT76), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n416_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n508_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT76), .B(new_n515_), .C1(new_n534_), .C2(new_n442_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n518_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n415_), .B(KEYINPUT36), .Z(new_n538_));
  NAND4_X1  g337(.A1(new_n537_), .A2(new_n528_), .A3(new_n519_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G1gat), .A2(G8gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT14), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(G1gat), .A2(G8gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .A4(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n551_), .B(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n564_), .A2(new_n566_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n560_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n511_), .A2(new_n559_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n510_), .A2(new_n482_), .A3(new_n474_), .A4(new_n558_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n559_), .A2(KEYINPUT12), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n534_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n574_), .A2(new_n583_), .A3(new_n576_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n578_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT5), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n578_), .B(new_n593_), .C1(new_n582_), .C2(new_n586_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(KEYINPUT13), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT13), .B1(new_n592_), .B2(new_n594_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n435_), .A2(new_n441_), .A3(new_n549_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n549_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n549_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n512_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n608_), .B2(new_n602_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  AND3_X1   g411(.A1(new_n605_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n600_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n605_), .A2(new_n609_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n605_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(KEYINPUT81), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n599_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n411_), .A2(new_n540_), .A3(new_n572_), .A4(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n367_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626_));
  INV_X1    g425(.A(new_n387_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n266_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n367_), .A2(new_n406_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n389_), .A2(KEYINPUT99), .A3(new_n392_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n392_), .B1(new_n389_), .B2(KEYINPUT99), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n403_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n634_), .B2(new_n266_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n410_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n635_), .A2(new_n636_), .B1(new_n345_), .B2(new_n385_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n622_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n598_), .B(KEYINPUT73), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n540_), .A2(KEYINPUT37), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT78), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n533_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT78), .B(new_n416_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n539_), .A2(KEYINPUT79), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n519_), .A2(new_n528_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT79), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .A4(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n640_), .B1(new_n648_), .B2(KEYINPUT37), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n571_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n638_), .A2(KEYINPUT104), .A3(new_n639_), .A4(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n411_), .A2(new_n621_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n639_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n367_), .A2(G1gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT105), .A3(new_n626_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT105), .B1(new_n657_), .B2(new_n626_), .ZN(new_n659_));
  OAI221_X1 g458(.A(new_n625_), .B1(new_n626_), .B2(new_n657_), .C1(new_n658_), .C2(new_n659_), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n343_), .A2(new_n344_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(G8gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n655_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT106), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n624_), .B2(new_n661_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT39), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(KEYINPUT40), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n624_), .B2(new_n636_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT41), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n638_), .A2(new_n639_), .A3(new_n650_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(G15gat), .A3(new_n636_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n624_), .B2(new_n408_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n408_), .A2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n674_), .B2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(new_n540_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n571_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n599_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n638_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n427_), .A3(new_n368_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n649_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n637_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n411_), .A2(new_n649_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n623_), .A2(new_n571_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n367_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n411_), .A2(new_n649_), .A3(new_n692_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n687_), .B1(new_n411_), .B2(new_n649_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n696_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n695_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(KEYINPUT44), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n699_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(KEYINPUT109), .A3(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT109), .B1(new_n707_), .B2(G29gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n686_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n705_), .A2(new_n704_), .A3(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n661_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n705_), .B2(KEYINPUT44), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n425_), .B1(new_n714_), .B2(new_n717_), .ZN(new_n718_));
  AND4_X1   g517(.A1(new_n425_), .A2(new_n638_), .A3(new_n715_), .A4(new_n683_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n711_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n720_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n716_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n722_), .B(KEYINPUT46), .C1(new_n425_), .C2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1329gat));
  OAI211_X1 g524(.A(G43gat), .B(new_n410_), .C1(new_n705_), .C2(KEYINPUT44), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G43gat), .B1(new_n685_), .B2(new_n410_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n727_), .A2(KEYINPUT47), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n727_), .B2(new_n728_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n685_), .A2(new_n418_), .A3(new_n266_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n408_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n714_), .B2(new_n734_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n736_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n637_), .A2(new_n621_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(new_n599_), .A3(new_n650_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n368_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT111), .Z(new_n742_));
  INV_X1    g541(.A(new_n639_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n621_), .A2(new_n571_), .ZN(new_n744_));
  AND4_X1   g543(.A1(new_n411_), .A2(new_n743_), .A3(new_n540_), .A4(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n368_), .A2(G57gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n745_), .B2(new_n715_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT48), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n740_), .A2(new_n748_), .A3(new_n715_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n740_), .A2(new_n753_), .A3(new_n410_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n745_), .A2(new_n410_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G71gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT113), .ZN(G1334gat));
  INV_X1    g559(.A(G78gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n745_), .B2(new_n266_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT50), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n740_), .A2(new_n761_), .A3(new_n266_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1335gat));
  NAND3_X1  g564(.A1(new_n599_), .A2(new_n622_), .A3(new_n571_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n367_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n639_), .A2(new_n682_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n739_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n368_), .A2(new_n460_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT114), .Z(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n768_), .B2(new_n661_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n771_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n461_), .A3(new_n715_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n768_), .B2(new_n636_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n410_), .A3(new_n479_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n266_), .A3(new_n444_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n492_), .B1(new_n767_), .B2(new_n266_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n783_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  XNOR2_X1  g591(.A(new_n744_), .B(KEYINPUT115), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n599_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n689_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT116), .B1(new_n795_), .B2(KEYINPUT54), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT54), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n689_), .A2(new_n794_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n601_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n608_), .A2(new_n602_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n802_), .B(new_n617_), .C1(new_n803_), .C2(new_n606_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n594_), .A2(new_n619_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n574_), .A2(new_n576_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT72), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n574_), .A2(new_n583_), .A3(new_n576_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n581_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n530_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n811_), .A2(new_n813_), .A3(KEYINPUT55), .A4(new_n580_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n574_), .B(new_n580_), .C1(new_n534_), .C2(new_n581_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n577_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n807_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n591_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n805_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI221_X1 g621(.A(new_n805_), .B1(KEYINPUT119), .B2(KEYINPUT58), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n649_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n594_), .A2(new_n621_), .A3(KEYINPUT117), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n594_), .B2(new_n621_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n592_), .A2(new_n594_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n619_), .A3(new_n804_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .A3(new_n540_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n681_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(KEYINPUT57), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n571_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n801_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n345_), .A2(new_n368_), .A3(new_n410_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n834_), .B2(KEYINPUT57), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(new_n830_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n817_), .A2(new_n591_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n827_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n843_), .B(new_n844_), .C1(new_n851_), .C2(new_n681_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n842_), .A2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n824_), .A2(new_n832_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT120), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n571_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n839_), .B1(new_n859_), .B2(new_n801_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n621_), .B(new_n841_), .C1(new_n860_), .C2(new_n838_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G113gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n801_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n840_), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n864_), .A2(G113gat), .A3(new_n622_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1340gat));
  OAI211_X1 g665(.A(new_n743_), .B(new_n841_), .C1(new_n860_), .C2(new_n838_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n860_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(G1341gat));
  OAI211_X1 g671(.A(new_n572_), .B(new_n841_), .C1(new_n860_), .C2(new_n838_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G127gat), .ZN(new_n874_));
  OR3_X1    g673(.A1(new_n864_), .A2(G127gat), .A3(new_n571_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1342gat));
  OAI211_X1 g675(.A(new_n649_), .B(new_n841_), .C1(new_n860_), .C2(new_n838_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G134gat), .ZN(new_n878_));
  OR3_X1    g677(.A1(new_n864_), .A2(G134gat), .A3(new_n540_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n410_), .A2(new_n408_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n661_), .A3(new_n368_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT121), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n863_), .A2(new_n621_), .A3(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n863_), .A2(new_n743_), .A3(new_n883_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g686(.A1(new_n863_), .A2(new_n572_), .A3(new_n883_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  INV_X1    g689(.A(G162gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n863_), .A2(new_n891_), .A3(new_n681_), .A4(new_n883_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n863_), .A2(new_n649_), .A3(new_n883_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1347gat));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n661_), .A2(new_n368_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n410_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n408_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n837_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n901_), .B2(new_n622_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n622_), .B(new_n899_), .C1(new_n801_), .C2(new_n836_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT122), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n904_), .A3(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n281_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n902_), .A2(new_n904_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(new_n266_), .B1(new_n859_), .B2(new_n801_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n743_), .A2(G176gat), .A3(new_n898_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n837_), .A2(new_n599_), .A3(new_n900_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n911_), .A2(new_n912_), .B1(new_n280_), .B2(new_n913_), .ZN(G1349gat));
  NOR3_X1   g713(.A1(new_n901_), .A2(new_n288_), .A3(new_n571_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n572_), .A3(new_n898_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n286_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n901_), .B2(new_n689_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n681_), .A2(new_n308_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT123), .Z(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n901_), .B2(new_n920_), .ZN(G1351gat));
  NAND2_X1  g720(.A1(new_n881_), .A2(new_n896_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n863_), .A2(G197gat), .A3(new_n621_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n863_), .A2(new_n621_), .A3(new_n923_), .ZN(new_n927_));
  INV_X1    g726(.A(G197gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n922_), .B1(new_n859_), .B2(new_n801_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n930_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n621_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n926_), .A2(new_n929_), .A3(new_n931_), .ZN(G1352gat));
  AND2_X1   g731(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n930_), .B(new_n743_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n863_), .A2(new_n923_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n639_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n937_), .B2(new_n934_), .ZN(G1353gat));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n930_), .B(new_n572_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n936_), .A2(new_n571_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n939_), .ZN(G1354gat));
  AND3_X1   g742(.A1(new_n930_), .A2(G218gat), .A3(new_n649_), .ZN(new_n944_));
  AOI211_X1 g743(.A(new_n540_), .B(new_n922_), .C1(new_n859_), .C2(new_n801_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G218gat), .B1(new_n945_), .B2(KEYINPUT126), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n936_), .B2(new_n540_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


