//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n208_), .A2(KEYINPUT24), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n204_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n209_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n206_), .A2(KEYINPUT22), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G169gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n221_), .A3(new_n207_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n210_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(KEYINPUT82), .A3(new_n210_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G15gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G71gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n231_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G127gat), .B(G134gat), .Z(new_n238_));
  XOR2_X1   g037(.A(G113gat), .B(G120gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n237_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT83), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT31), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  AND2_X1   g049(.A1(G197gat), .A2(G204gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254_));
  AOI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G211gat), .B(G218gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT21), .B2(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n223_), .A2(KEYINPUT94), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n213_), .A2(new_n226_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n222_), .B2(new_n210_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n204_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n216_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n261_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n259_), .A2(KEYINPUT21), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n259_), .B2(new_n255_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n218_), .A3(new_n229_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(KEYINPUT20), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT19), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G8gat), .B(G36gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n268_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n214_), .B1(KEYINPUT24), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n265_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n227_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n272_), .B(new_n285_), .C1(new_n262_), .C2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n230_), .A2(new_n261_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n276_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT20), .A4(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n277_), .A2(new_n283_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT20), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n276_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(KEYINPUT99), .A3(new_n276_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n296_), .B(new_n297_), .C1(new_n276_), .C2(new_n274_), .ZN(new_n298_));
  AOI211_X1 g097(.A(new_n249_), .B(new_n292_), .C1(new_n298_), .C2(new_n282_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n283_), .B1(new_n277_), .B2(new_n291_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n292_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT27), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT96), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(G155gat), .A3(G162gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G141gat), .ZN(new_n312_));
  INV_X1    g111(.A(G148gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT84), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n314_), .A2(new_n316_), .B1(G141gat), .B2(G148gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT85), .A3(new_n311_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n318_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  OAI22_X1  g127(.A1(KEYINPUT86), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n310_), .A2(new_n306_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n321_), .A2(new_n323_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n240_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n331_), .ZN(new_n334_));
  AND4_X1   g133(.A1(KEYINPUT85), .A2(new_n311_), .A3(new_n318_), .A4(new_n317_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT85), .B1(new_n322_), .B2(new_n311_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n241_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n338_), .A3(KEYINPUT4), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n240_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n305_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n333_), .A2(new_n338_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(new_n304_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n299_), .A2(new_n302_), .A3(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G22gat), .B(G50gat), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n332_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n359_), .A2(new_n360_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n357_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT88), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n261_), .B(new_n373_), .C1(new_n332_), .C2(new_n358_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n272_), .B1(new_n337_), .B2(KEYINPUT29), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n370_), .B(KEYINPUT90), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n374_), .B(KEYINPUT91), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n321_), .A2(new_n323_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n358_), .B1(new_n380_), .B2(new_n334_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n381_), .B2(new_n272_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT91), .B1(new_n382_), .B2(new_n374_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n368_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  INV_X1    g184(.A(new_n368_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n374_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n376_), .B1(new_n388_), .B2(new_n261_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n384_), .A2(new_n385_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT92), .B(new_n368_), .C1(new_n378_), .C2(new_n383_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n367_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n386_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n368_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n367_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT93), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n367_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n386_), .B1(new_n400_), .B2(new_n377_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n401_), .B2(KEYINPUT92), .ZN(new_n402_));
  INV_X1    g201(.A(new_n392_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n398_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n396_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n355_), .A2(new_n397_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n353_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT33), .B(new_n350_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n339_), .A2(new_n340_), .A3(new_n305_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n343_), .A2(new_n304_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n351_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n301_), .A2(new_n410_), .A3(new_n411_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n298_), .A2(KEYINPUT32), .A3(new_n283_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n274_), .A2(new_n276_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n291_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n283_), .A2(KEYINPUT32), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n352_), .A2(new_n353_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n415_), .A2(KEYINPUT98), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n412_), .A2(new_n413_), .A3(new_n351_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n292_), .A2(new_n423_), .A3(new_n300_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT98), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n397_), .A2(new_n407_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n408_), .B1(new_n427_), .B2(KEYINPUT100), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n415_), .A2(KEYINPUT98), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n421_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n384_), .A2(new_n385_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n433_));
  AOI211_X1 g232(.A(KEYINPUT93), .B(new_n396_), .C1(new_n433_), .C2(new_n398_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n406_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT100), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n248_), .B1(new_n428_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT101), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT101), .B(new_n248_), .C1(new_n428_), .C2(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n397_), .A2(new_n407_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n299_), .A2(new_n302_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n445_), .A2(new_n248_), .A3(new_n354_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n441_), .A2(new_n442_), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G169gat), .B(G197gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT77), .B(G15gat), .ZN(new_n453_));
  INV_X1    g252(.A(G22gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n460_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n466_), .A2(KEYINPUT80), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(KEYINPUT80), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n462_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n465_), .B(KEYINPUT15), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n465_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n452_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n467_), .A2(new_n468_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n479_), .B(new_n451_), .C1(new_n470_), .C2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n448_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G232gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT34), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(KEYINPUT75), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT6), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  OR3_X1    g291(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT8), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  INV_X1    g300(.A(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n495_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n496_), .B1(new_n495_), .B2(KEYINPUT9), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n491_), .B(new_n503_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n500_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n512_), .A2(new_n513_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n517_), .A2(new_n465_), .B1(new_n487_), .B2(new_n486_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT69), .B1(new_n515_), .B2(new_n516_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n516_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n514_), .A4(new_n500_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n472_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n489_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n488_), .A2(KEYINPUT75), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n523_), .A3(KEYINPUT75), .A4(new_n488_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT36), .Z(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(KEYINPUT36), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT76), .B1(new_n528_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT76), .ZN(new_n537_));
  INV_X1    g336(.A(new_n535_), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n537_), .B(new_n538_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n534_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n534_), .B(KEYINPUT37), .C1(new_n536_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT11), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(new_n546_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n471_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT78), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n557_), .B(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n555_), .A2(KEYINPUT17), .A3(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n544_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT79), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n552_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n520_), .A2(new_n514_), .A3(new_n500_), .A4(new_n551_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n517_), .A2(KEYINPUT68), .A3(new_n551_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n519_), .A2(new_n522_), .A3(KEYINPUT12), .A4(new_n552_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n569_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n571_), .A2(KEYINPUT70), .A3(new_n573_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT70), .B1(new_n571_), .B2(new_n573_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n576_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n576_), .B(new_n590_), .C1(new_n580_), .C2(new_n583_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT73), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(KEYINPUT73), .A3(new_n594_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT13), .B1(new_n596_), .B2(new_n597_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT74), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n483_), .A2(new_n568_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n456_), .A3(new_n354_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n602_), .A2(new_n482_), .A3(new_n604_), .A4(new_n565_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT102), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n540_), .B(KEYINPUT103), .Z(new_n612_));
  AOI21_X1  g411(.A(new_n446_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(new_n442_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n354_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n607_), .A2(new_n608_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(new_n444_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n606_), .A2(new_n457_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n615_), .B2(new_n444_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1325gat));
  INV_X1    g426(.A(new_n248_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n628_), .A3(new_n614_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(G15gat), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(new_n634_), .A3(new_n632_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n606_), .A2(new_n233_), .A3(new_n628_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(G1326gat));
  NOR2_X1   g438(.A1(new_n434_), .A2(new_n435_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n606_), .A2(new_n454_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n615_), .B2(new_n443_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n641_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT106), .ZN(G1327gat));
  INV_X1    g445(.A(new_n482_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n613_), .B2(new_n442_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n540_), .A2(new_n565_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n605_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n354_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n605_), .A2(new_n647_), .A3(new_n565_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n544_), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT43), .B(new_n656_), .C1(new_n613_), .C2(new_n442_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n448_), .B2(new_n544_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n655_), .B(KEYINPUT44), .C1(new_n657_), .C2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(G29gat), .A3(new_n354_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n655_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n654_), .B1(new_n661_), .B2(new_n664_), .ZN(G1328gat));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n620_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n436_), .A2(new_n437_), .B1(new_n640_), .B2(new_n355_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n427_), .A2(KEYINPUT100), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n628_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n447_), .B1(new_n669_), .B2(KEYINPUT101), .ZN(new_n670_));
  INV_X1    g469(.A(new_n442_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n544_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT43), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n448_), .A2(new_n658_), .A3(new_n544_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n675_), .B2(new_n655_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G36gat), .B1(new_n666_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n444_), .A2(G36gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n653_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n653_), .A2(new_n682_), .A3(new_n679_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n677_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n660_), .A2(G43gat), .A3(new_n628_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n652_), .A2(new_n248_), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n688_), .A2(new_n676_), .B1(G43gat), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n653_), .A2(new_n692_), .A3(new_n640_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n664_), .A2(new_n640_), .A3(new_n660_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(KEYINPUT108), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n664_), .A2(new_n696_), .A3(new_n640_), .A4(new_n660_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT109), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n660_), .A2(new_n640_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT108), .B1(new_n699_), .B2(new_n676_), .ZN(new_n700_));
  AND4_X1   g499(.A1(KEYINPUT109), .A2(new_n700_), .A3(G50gat), .A4(new_n697_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n693_), .B1(new_n698_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n605_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n568_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n482_), .B1(new_n613_), .B2(new_n442_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n354_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n565_), .A2(new_n647_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n703_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n614_), .A2(new_n710_), .A3(G57gat), .A4(new_n354_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n708_), .A2(new_n712_), .A3(new_n713_), .ZN(G1332gat));
  NAND2_X1  g513(.A1(new_n614_), .A2(new_n710_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G64gat), .B1(new_n715_), .B2(new_n444_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT48), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n444_), .A2(G64gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n706_), .B2(new_n718_), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n715_), .B2(new_n248_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT49), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n248_), .A2(G71gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n706_), .B2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n715_), .B2(new_n443_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n443_), .A2(G78gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n706_), .B2(new_n726_), .ZN(G1335gat));
  AND3_X1   g526(.A1(new_n705_), .A2(new_n605_), .A3(new_n649_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n354_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n605_), .A2(new_n647_), .A3(new_n566_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n675_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n354_), .A2(G85gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n730_), .B1(new_n734_), .B2(new_n736_), .ZN(G1336gat));
  INV_X1    g536(.A(G92gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n738_), .A3(new_n620_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n734_), .A2(new_n620_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n738_), .ZN(G1337gat));
  NAND3_X1  g541(.A1(new_n728_), .A2(new_n628_), .A3(new_n501_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(KEYINPUT114), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n734_), .A2(new_n628_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G99gat), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n744_), .A2(KEYINPUT114), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n728_), .A2(new_n502_), .A3(new_n640_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n675_), .A2(new_n733_), .A3(new_n640_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G106gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G106gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n647_), .B(new_n565_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n544_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n600_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n709_), .B1(new_n763_), .B2(new_n598_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n656_), .A2(new_n764_), .A3(new_n759_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n758_), .B1(new_n762_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n470_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n469_), .A2(new_n767_), .A3(new_n473_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n452_), .C1(new_n767_), .C2(new_n480_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n481_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n594_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n571_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n574_), .B1(new_n580_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n776_));
  OR3_X1    g575(.A1(new_n580_), .A2(new_n583_), .A3(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT118), .B(new_n574_), .C1(new_n580_), .C2(new_n772_), .ZN(new_n778_));
  AND2_X1   g577(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n779_));
  OAI22_X1  g578(.A1(new_n580_), .A2(new_n583_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n775_), .A2(new_n777_), .A3(new_n778_), .A4(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n591_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT58), .B(new_n771_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT120), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n591_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n591_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT58), .A4(new_n771_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n771_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n785_), .A2(new_n792_), .A3(new_n795_), .A4(new_n544_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n482_), .A2(new_n594_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n482_), .A2(KEYINPUT116), .A3(new_n594_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n596_), .A2(new_n597_), .A3(new_n770_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n540_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n799_), .B(new_n800_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n803_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n540_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n796_), .A2(new_n807_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n766_), .B1(new_n811_), .B2(new_n566_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n248_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n445_), .A2(new_n616_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n482_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n647_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n818_), .B1(new_n821_), .B2(new_n817_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n703_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n816_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n703_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n816_), .A2(new_n828_), .A3(new_n565_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n566_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n816_), .B2(new_n612_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n819_), .A2(new_n820_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT121), .B(G134gat), .Z(new_n834_));
  NOR2_X1   g633(.A1(new_n656_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n811_), .A2(new_n566_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n766_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n628_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(new_n640_), .A3(new_n354_), .A4(new_n444_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n647_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n312_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n703_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n313_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n840_), .A2(new_n566_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  OAI21_X1  g646(.A(G162gat), .B1(new_n840_), .B2(new_n656_), .ZN(new_n848_));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n612_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n840_), .B2(new_n850_), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n444_), .A2(new_n354_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n640_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n813_), .A2(new_n482_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT122), .B1(new_n855_), .B2(G169gat), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n219_), .A2(new_n221_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n860_), .B(new_n861_), .C1(new_n862_), .C2(new_n855_), .ZN(G1348gat));
  NAND2_X1  g662(.A1(new_n813_), .A2(new_n854_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n703_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT123), .B(G176gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1349gat));
  NAND3_X1  g666(.A1(new_n813_), .A2(new_n565_), .A3(new_n854_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G183gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n202_), .B1(KEYINPUT124), .B2(G183gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n868_), .B2(new_n871_), .ZN(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n864_), .B2(new_n656_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n612_), .A2(new_n203_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n864_), .B2(new_n874_), .ZN(G1351gat));
  NOR2_X1   g674(.A1(new_n853_), .A2(new_n443_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n809_), .B2(new_n540_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n540_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n806_), .B(new_n878_), .C1(new_n808_), .C2(new_n803_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n565_), .B1(new_n880_), .B2(new_n796_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n248_), .B(new_n876_), .C1(new_n881_), .C2(new_n766_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT125), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n839_), .A2(new_n884_), .A3(new_n876_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n482_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT126), .B(G204gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n605_), .ZN(new_n891_));
  MUX2_X1   g690(.A(new_n889_), .B(new_n890_), .S(new_n891_), .Z(G1353gat));
  OR2_X1    g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND4_X1   g693(.A1(new_n565_), .A2(new_n886_), .A3(new_n893_), .A4(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n886_), .B2(new_n565_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n884_), .B1(new_n839_), .B2(new_n876_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n876_), .ZN(new_n900_));
  NOR4_X1   g699(.A1(new_n812_), .A2(KEYINPUT125), .A3(new_n628_), .A4(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n898_), .B(new_n612_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n656_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n902_), .B(new_n903_), .C1(new_n904_), .C2(new_n898_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n544_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G218gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n903_), .B1(new_n908_), .B2(new_n902_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n906_), .A2(new_n909_), .ZN(G1355gat));
endmodule


