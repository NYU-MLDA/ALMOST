//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT66), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n211_), .A2(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n207_), .A2(KEYINPUT66), .ZN(new_n218_));
  OAI211_X1 g017(.A(KEYINPUT8), .B(new_n202_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n207_), .A3(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n202_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n215_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(G92gat), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n224_), .A2(new_n226_), .A3(new_n230_), .A4(new_n207_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n219_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G57gat), .B(G64gat), .Z(new_n233_));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT67), .B(G71gat), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(G78gat), .ZN(new_n239_));
  AND4_X1   g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n235_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n232_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT12), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n232_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G176gat), .B(G204gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(G120gat), .B(G148gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n249_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT13), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT13), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(KEYINPUT69), .A3(new_n264_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G113gat), .B(G120gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273_));
  INV_X1    g072(.A(G155gat), .ZN(new_n274_));
  INV_X1    g073(.A(G162gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT91), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT2), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(KEYINPUT90), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n286_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n279_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n278_), .A2(KEYINPUT1), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(G155gat), .A3(G162gat), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n276_), .A2(new_n290_), .A3(new_n292_), .A4(new_n277_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n283_), .A2(new_n284_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n272_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT2), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n280_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n300_), .A2(new_n302_), .A3(new_n287_), .A4(new_n285_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n279_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n271_), .B(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n297_), .A2(KEYINPUT4), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G1gat), .B(G29gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G85gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT0), .B(G57gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  AOI21_X1  g120(.A(new_n316_), .B1(new_n297_), .B2(new_n309_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n315_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT86), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n330_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G71gat), .B(G99gat), .Z(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G15gat), .B(G43gat), .Z(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n336_), .A3(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT87), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT31), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n345_), .A2(KEYINPUT87), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n345_), .B2(KEYINPUT87), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  NOR4_X1   g152(.A1(new_n343_), .A2(new_n344_), .A3(new_n353_), .A4(KEYINPUT31), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT88), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n361_));
  OAI22_X1  g160(.A1(new_n358_), .A2(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G169gat), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n366_), .A3(new_n371_), .A4(KEYINPUT81), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT82), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(KEYINPUT82), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n374_), .A2(new_n375_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n380_), .A2(new_n381_), .ZN(new_n386_));
  INV_X1    g185(.A(G183gat), .ZN(new_n387_));
  INV_X1    g186(.A(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n365_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G169gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n367_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n368_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n395_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT30), .B1(new_n385_), .B2(new_n399_), .ZN(new_n400_));
  OR3_X1    g199(.A1(new_n385_), .A2(new_n399_), .A3(KEYINPUT30), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n357_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n307_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n357_), .A2(new_n401_), .A3(new_n272_), .A4(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n356_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n351_), .A2(new_n355_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n329_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n414_));
  INV_X1    g213(.A(G204gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G197gat), .ZN(new_n416_));
  INV_X1    g215(.A(G197gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G204gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G211gat), .B(G218gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n421_), .B(new_n420_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(G228gat), .B(G233gat), .C1(new_n414_), .C2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G22gat), .B(G50gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n305_), .A2(new_n308_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(KEYINPUT29), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n305_), .A2(new_n434_), .A3(new_n308_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(KEYINPUT29), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n427_), .A2(new_n439_), .A3(new_n428_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT94), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n427_), .A2(new_n439_), .A3(new_n428_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n430_), .B(new_n437_), .C1(new_n441_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT94), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n437_), .B1(new_n450_), .B2(new_n430_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n412_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n430_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n437_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(new_n411_), .A3(new_n446_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT27), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n427_), .A2(new_n428_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n385_), .B2(new_n399_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n359_), .A2(new_n358_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n360_), .A2(new_n361_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT97), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n466_), .A2(new_n467_), .B1(new_n382_), .B2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n377_), .A2(new_n380_), .A3(KEYINPUT97), .A4(new_n381_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n369_), .A2(KEYINPUT24), .A3(new_n370_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n368_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n469_), .A2(new_n472_), .B1(new_n390_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n465_), .B1(new_n478_), .B2(new_n429_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n461_), .A2(new_n464_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n463_), .B(KEYINPUT96), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n374_), .A2(new_n375_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n383_), .A2(new_n384_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n429_), .A3(new_n398_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n390_), .A2(new_n477_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n382_), .A2(new_n468_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n487_), .A2(new_n471_), .A3(new_n362_), .A4(new_n470_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n465_), .B1(new_n489_), .B2(new_n460_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n481_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT18), .B(G64gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n480_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n481_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n385_), .A2(new_n399_), .A3(new_n460_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n478_), .B2(new_n429_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n461_), .A2(new_n464_), .A3(new_n479_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n496_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n459_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n489_), .B2(new_n460_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT99), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n479_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n510_), .A3(new_n461_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n500_), .A2(new_n501_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n511_), .A2(new_n463_), .B1(new_n512_), .B2(new_n481_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT27), .B(new_n506_), .C1(new_n513_), .C2(new_n496_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n458_), .A2(new_n505_), .A3(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n408_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n406_), .A2(new_n407_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n498_), .A2(new_n504_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n297_), .A2(new_n316_), .A3(new_n309_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n321_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n310_), .A2(new_n315_), .A3(new_n313_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n327_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(KEYINPUT33), .B(new_n325_), .C1(new_n326_), .C2(new_n322_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT98), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n317_), .A2(new_n323_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT33), .A4(new_n325_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n518_), .A2(new_n524_), .A3(new_n526_), .A4(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n496_), .A2(KEYINPUT32), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n502_), .A2(new_n531_), .A3(new_n503_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n328_), .B(new_n532_), .C1(new_n513_), .C2(new_n531_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n457_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n328_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n535_), .A2(new_n505_), .A3(new_n514_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n517_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n516_), .B1(new_n537_), .B2(KEYINPUT100), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n517_), .C1(new_n534_), .C2(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT74), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G15gat), .ZN(new_n545_));
  INV_X1    g344(.A(G22gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G15gat), .A2(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G1gat), .A2(G8gat), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n547_), .A2(new_n548_), .B1(KEYINPUT14), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n544_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G43gat), .B(G50gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n551_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n551_), .A2(new_n556_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT15), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n556_), .B(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n565_), .B2(new_n551_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n558_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT78), .B(G169gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G197gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n568_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT79), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n269_), .A2(new_n541_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n242_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(new_n551_), .Z(new_n579_));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G211gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT16), .B(G183gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT76), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  INV_X1    g388(.A(new_n579_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(KEYINPUT76), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n588_), .B2(new_n592_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n565_), .A2(new_n232_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n556_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n219_), .A2(new_n223_), .A3(new_n598_), .A4(new_n231_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(KEYINPUT71), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT35), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n565_), .A2(new_n232_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  INV_X1    g412(.A(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n605_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n597_), .A2(new_n614_), .A3(new_n599_), .A4(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n609_), .A2(new_n610_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n613_), .B(KEYINPUT36), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n609_), .A2(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT73), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT73), .B1(new_n609_), .B2(new_n616_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n617_), .B(new_n618_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n620_), .A2(new_n619_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n617_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT37), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT72), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n596_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n576_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G1gat), .A3(new_n329_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT101), .Z(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n269_), .A2(new_n575_), .A3(new_n595_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT102), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n622_), .A2(new_n623_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n617_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT103), .Z(new_n644_));
  AND2_X1   g443(.A1(new_n541_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n329_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n638_), .A2(new_n639_), .A3(new_n647_), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n514_), .A2(new_n505_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n634_), .A2(G8gat), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G8gat), .B1(new_n646_), .B2(new_n649_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g454(.A(new_n634_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n407_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n351_), .A2(new_n355_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n545_), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G15gat), .B1(new_n646_), .B2(new_n517_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n546_), .A3(new_n457_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G22gat), .B1(new_n646_), .B2(new_n458_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  XOR2_X1   g469(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n671_));
  NAND4_X1  g470(.A1(new_n267_), .A2(new_n596_), .A3(new_n575_), .A4(new_n268_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n629_), .A2(new_n631_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(KEYINPUT104), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n676_), .B(new_n673_), .C1(new_n675_), .C2(KEYINPUT104), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT106), .B(new_n672_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n659_), .A2(new_n649_), .A3(new_n329_), .A4(new_n458_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n497_), .B1(new_n480_), .B2(new_n491_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n327_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n523_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(new_n506_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n529_), .A2(new_n526_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n533_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n458_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n535_), .A2(new_n505_), .A3(new_n514_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n659_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n692_), .B2(new_n539_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n540_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n632_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n695_), .B2(KEYINPUT105), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT105), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n680_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n672_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n682_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n671_), .B1(new_n681_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT108), .B(new_n671_), .C1(new_n681_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n672_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(KEYINPUT44), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n707_), .A2(new_n699_), .A3(KEYINPUT44), .A4(new_n700_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n328_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n706_), .A2(KEYINPUT110), .A3(new_n328_), .A4(new_n713_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(G29gat), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n643_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n596_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n576_), .A2(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n329_), .A2(G29gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n649_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n713_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  INV_X1    g527(.A(new_n722_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n649_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n725_), .A3(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT45), .Z(new_n732_));
  OR3_X1    g531(.A1(new_n727_), .A2(new_n728_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n728_), .B1(new_n727_), .B2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n722_), .B2(new_n517_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n517_), .A2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT111), .B(new_n739_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741_));
  INV_X1    g540(.A(new_n739_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n706_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n737_), .C1(new_n740_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1330gat));
  AOI21_X1  g547(.A(G50gat), .B1(new_n729_), .B2(new_n457_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n706_), .A2(G50gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n458_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n269_), .A2(new_n575_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n541_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n633_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n328_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n644_), .A3(new_n595_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n329_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(G57gat), .B2(new_n759_), .ZN(G1332gat));
  OR3_X1    g559(.A1(new_n755_), .A2(G64gat), .A3(new_n649_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G64gat), .B1(new_n758_), .B2(new_n649_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1333gat));
  OR3_X1    g567(.A1(new_n755_), .A2(G71gat), .A3(new_n517_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G71gat), .B1(new_n758_), .B2(new_n517_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n770_), .A2(KEYINPUT49), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n770_), .A2(KEYINPUT49), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n758_), .B2(new_n458_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n458_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n755_), .B2(new_n779_), .ZN(G1335gat));
  NAND2_X1  g579(.A1(new_n754_), .A2(new_n721_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n328_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n699_), .A2(new_n596_), .A3(new_n753_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n229_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n329_), .B1(new_n785_), .B2(new_n227_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(G1336gat));
  AOI21_X1  g586(.A(G92gat), .B1(new_n782_), .B2(new_n730_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n649_), .A2(new_n493_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT114), .ZN(G1337gat));
  AOI21_X1  g590(.A(new_n214_), .B1(new_n784_), .B2(new_n659_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT115), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n782_), .A2(new_n225_), .A3(new_n659_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g595(.A1(new_n784_), .A2(new_n457_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G106gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT116), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT52), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n782_), .A2(new_n215_), .A3(new_n457_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n806_), .B(new_n808_), .ZN(G1339gat));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n517_), .A2(new_n515_), .A3(new_n329_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT55), .B1(new_n247_), .B2(new_n248_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n816_), .B(new_n250_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n247_), .A2(new_n248_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n815_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n813_), .B(new_n814_), .C1(new_n819_), .C2(new_n257_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n815_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n817_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n818_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n258_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n258_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n813_), .B1(new_n827_), .B2(new_n814_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n575_), .B(new_n260_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n568_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n557_), .A2(new_n558_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n572_), .B1(new_n566_), .B2(new_n559_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n830_), .A2(new_n572_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n261_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n643_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n835_), .A2(new_n643_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n825_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n260_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n827_), .A2(new_n814_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n842_), .A3(new_n825_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n833_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n833_), .A4(new_n847_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n632_), .A3(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n839_), .A2(new_n841_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n596_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n596_), .B2(new_n575_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n573_), .B(KEYINPUT79), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT118), .A3(new_n595_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n856_), .A2(new_n265_), .A3(new_n674_), .A4(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT54), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT59), .B(new_n812_), .C1(new_n854_), .C2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n840_), .B1(new_n835_), .B2(new_n643_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n719_), .B(new_n838_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n595_), .B1(new_n864_), .B2(new_n852_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n860_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n854_), .A2(new_n868_), .A3(new_n860_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n869_), .A3(new_n811_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n810_), .B(new_n861_), .C1(new_n870_), .C2(KEYINPUT59), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n867_), .A2(new_n869_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n575_), .A3(new_n811_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n871_), .A2(new_n575_), .B1(new_n810_), .B2(new_n873_), .ZN(G1340gat));
  AOI211_X1 g673(.A(new_n269_), .B(new_n861_), .C1(new_n870_), .C2(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(KEYINPUT60), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n269_), .B2(KEYINPUT60), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n811_), .A3(new_n878_), .ZN(new_n879_));
  OAI22_X1  g678(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1341gat));
  NOR2_X1   g679(.A1(KEYINPUT123), .A2(G127gat), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n881_), .B(new_n861_), .C1(new_n870_), .C2(KEYINPUT59), .ZN(new_n882_));
  OAI21_X1  g681(.A(G127gat), .B1(new_n596_), .B2(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n872_), .A2(new_n595_), .A3(new_n811_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n882_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1342gat));
  XOR2_X1   g685(.A(KEYINPUT124), .B(G134gat), .Z(new_n887_));
  AOI211_X1 g686(.A(new_n887_), .B(new_n861_), .C1(new_n870_), .C2(KEYINPUT59), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n644_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n872_), .A2(new_n890_), .A3(new_n811_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n888_), .A2(new_n632_), .B1(new_n889_), .B2(new_n891_), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n730_), .A2(new_n458_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n872_), .A2(new_n328_), .A3(new_n517_), .A4(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894_), .B2(new_n857_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n867_), .A2(new_n869_), .A3(new_n328_), .A4(new_n517_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n896_), .A2(new_n458_), .A3(new_n730_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n283_), .A3(new_n575_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1344gat));
  OAI21_X1  g698(.A(G148gat), .B1(new_n894_), .B2(new_n269_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n269_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n284_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1345gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n897_), .A2(new_n595_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n897_), .B2(new_n595_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1346gat));
  NOR3_X1   g706(.A1(new_n894_), .A2(new_n275_), .A3(new_n674_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G162gat), .B1(new_n897_), .B2(new_n890_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n854_), .A2(new_n860_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n408_), .A2(new_n649_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n458_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT125), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n911_), .A2(new_n915_), .A3(new_n458_), .A4(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(new_n476_), .A3(new_n575_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n913_), .A2(new_n857_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n919_), .A2(new_n920_), .A3(G169gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(G169gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n918_), .B1(new_n921_), .B2(new_n922_), .ZN(G1348gat));
  AOI21_X1  g722(.A(G176gat), .B1(new_n917_), .B2(new_n901_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n867_), .A2(new_n869_), .A3(new_n458_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n867_), .A2(new_n869_), .A3(KEYINPUT126), .A4(new_n458_), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n368_), .B(new_n269_), .C1(new_n927_), .C2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n924_), .B1(new_n929_), .B2(new_n912_), .ZN(G1349gat));
  AOI211_X1 g729(.A(new_n466_), .B(new_n596_), .C1(new_n914_), .C2(new_n916_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n928_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(new_n595_), .A3(new_n912_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(new_n387_), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n917_), .A2(new_n890_), .A3(new_n467_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n674_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n388_), .ZN(G1351gat));
  NAND4_X1  g736(.A1(new_n867_), .A2(new_n869_), .A3(new_n535_), .A4(new_n517_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n938_), .A2(new_n649_), .A3(new_n857_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT127), .B(G197gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1352gat));
  NOR2_X1   g740(.A1(new_n938_), .A2(new_n649_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n901_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g743(.A(KEYINPUT63), .B(G211gat), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n938_), .A2(new_n649_), .A3(new_n596_), .A4(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n595_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n942_), .B2(new_n890_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n942_), .A2(G218gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n632_), .B2(new_n951_), .ZN(G1355gat));
endmodule


