//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT26), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G190gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT82), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT81), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n215_), .A2(new_n224_), .A3(KEYINPUT24), .A4(new_n216_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT83), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT23), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n226_), .A2(KEYINPUT23), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n223_), .B(new_n225_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n229_), .ZN(new_n235_));
  AOI211_X1 g034(.A(new_n233_), .B(new_n234_), .C1(new_n235_), .C2(KEYINPUT23), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT22), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n240_), .A3(new_n214_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n216_), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n222_), .A2(new_n232_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  INV_X1    g043(.A(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G15gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n247_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT85), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n259_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n258_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT85), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT86), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT31), .Z(new_n266_));
  NAND3_X1  g065(.A1(new_n254_), .A2(new_n255_), .A3(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n255_), .A2(new_n266_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT97), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OR3_X1    g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT19), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT94), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n286_), .B(new_n287_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n284_), .A2(new_n285_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n289_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n243_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n239_), .A2(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n213_), .A2(KEYINPUT22), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT95), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT95), .B1(new_n299_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n214_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n230_), .A2(new_n231_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n303_), .B(new_n216_), .C1(new_n304_), .C2(new_n233_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n234_), .B1(new_n235_), .B2(KEYINPUT23), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n306_), .A2(new_n210_), .A3(new_n217_), .A4(new_n223_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n305_), .A2(new_n307_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n283_), .B1(new_n298_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n243_), .A2(new_n297_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n305_), .A2(new_n296_), .A3(new_n292_), .A4(new_n307_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT20), .A4(new_n282_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n280_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G148gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(KEYINPUT3), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT89), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n318_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n324_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n328_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT88), .B1(new_n328_), .B2(KEYINPUT1), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G141gat), .B(G148gat), .Z(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n261_), .A2(new_n262_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n332_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n332_), .A2(new_n339_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT4), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n264_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G85gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n332_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n345_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n350_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n350_), .B2(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n313_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT20), .ZN(new_n361_));
  INV_X1    g160(.A(new_n282_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n298_), .A2(new_n308_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n283_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n363_), .A2(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(KEYINPUT100), .A3(new_n362_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n280_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT101), .B1(new_n360_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n350_), .A2(new_n357_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n354_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n350_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(new_n364_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n365_), .A2(new_n366_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n368_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n280_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT101), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n375_), .A2(new_n380_), .A3(new_n381_), .A4(new_n313_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n347_), .A2(new_n355_), .A3(new_n345_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n343_), .A2(new_n349_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT99), .B1(new_n384_), .B2(new_n344_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n386_), .B(new_n345_), .C1(new_n343_), .C2(new_n349_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n354_), .B(new_n383_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT98), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT33), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT4), .B1(new_n346_), .B2(new_n264_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n347_), .A2(new_n355_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT4), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n356_), .B1(new_n393_), .B2(new_n345_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n390_), .B1(new_n394_), .B2(new_n354_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n309_), .A2(new_n279_), .A3(new_n312_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n279_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n390_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n359_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n388_), .A2(new_n395_), .A3(new_n398_), .A4(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n370_), .A2(new_n382_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n346_), .A2(KEYINPUT29), .ZN(new_n403_));
  INV_X1    g202(.A(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(G228gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(G228gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n297_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n408_), .B(new_n409_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n292_), .A2(new_n296_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n346_), .A2(KEYINPUT29), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT28), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n422_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n411_), .A2(new_n416_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n417_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n419_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n428_), .A2(new_n425_), .A3(KEYINPUT93), .A4(new_n419_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n402_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n309_), .A2(new_n279_), .A3(new_n312_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT27), .ZN(new_n435_));
  INV_X1    g234(.A(new_n279_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n378_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n309_), .A2(new_n312_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n434_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT102), .A3(new_n438_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n437_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n432_), .A2(new_n375_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n269_), .B1(new_n433_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n375_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n267_), .A2(new_n450_), .A3(new_n268_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n378_), .A2(new_n436_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n435_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT102), .B1(new_n444_), .B2(new_n438_), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n440_), .B(KEYINPUT27), .C1(new_n443_), .C2(new_n434_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n432_), .B(new_n454_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT103), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n446_), .A2(KEYINPUT103), .A3(new_n432_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n451_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n449_), .A2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT65), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(KEYINPUT65), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n463_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT10), .B(G99gat), .Z(new_n473_));
  INV_X1    g272(.A(G106gat), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n469_), .A2(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT9), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(KEYINPUT64), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(KEYINPUT64), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n479_), .B(new_n478_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n475_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n475_), .B2(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n474_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G85gat), .B(G92gat), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n496_), .A2(KEYINPUT8), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n493_), .A2(new_n494_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n470_), .A2(new_n471_), .A3(new_n463_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n463_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n504_), .B2(new_n497_), .ZN(new_n505_));
  OAI22_X1  g304(.A1(new_n489_), .A2(new_n490_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n509_));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n509_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(KEYINPUT12), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n475_), .A2(new_n487_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT66), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n475_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT8), .B1(new_n496_), .B2(new_n498_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n504_), .A2(new_n500_), .A3(new_n497_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n522_), .A3(new_n513_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n515_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n506_), .A2(new_n514_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n506_), .C2(new_n514_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n524_), .B(new_n525_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n523_), .A3(KEYINPUT67), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n506_), .A2(KEYINPUT67), .A3(new_n514_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(G230gat), .A4(G233gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G176gat), .B(G204gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT70), .ZN(new_n537_));
  XOR2_X1   g336(.A(G120gat), .B(G148gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT13), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT13), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549_));
  XOR2_X1   g348(.A(G29gat), .B(G36gat), .Z(new_n550_));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT71), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n549_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n554_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n555_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT15), .A3(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565_));
  INV_X1    g364(.A(G1gat), .ZN(new_n566_));
  INV_X1    g365(.A(G8gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G8gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n556_), .A2(new_n557_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n573_), .B(new_n571_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT80), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G113gat), .B(G141gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G169gat), .B(G197gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n582_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n548_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n462_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT75), .ZN(new_n590_));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n558_), .A2(new_n563_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n522_), .B2(new_n519_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n506_), .A2(new_n573_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n564_), .A2(new_n506_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n599_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n605_), .B2(new_n599_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n595_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT35), .B(new_n601_), .C1(new_n597_), .C2(KEYINPUT72), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n603_), .B1(new_n506_), .B2(new_n573_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n595_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n607_), .A3(new_n615_), .A4(new_n609_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n611_), .A2(KEYINPUT37), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT37), .B1(new_n611_), .B2(new_n616_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT79), .ZN(new_n622_));
  XOR2_X1   g421(.A(G183gat), .B(G211gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT77), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n513_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n571_), .B(KEYINPUT76), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n632_), .A2(new_n634_), .A3(new_n626_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n620_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n588_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT104), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n566_), .A3(new_n375_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n611_), .A2(new_n616_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n462_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n636_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n548_), .A4(new_n586_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n450_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n640_), .A2(new_n641_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  OAI21_X1  g449(.A(G8gat), .B1(new_n647_), .B2(new_n446_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT39), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n446_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n639_), .A2(new_n567_), .A3(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n654_), .B(new_n656_), .C1(KEYINPUT39), .C2(new_n653_), .ZN(new_n657_));
  XOR2_X1   g456(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  NAND3_X1  g458(.A1(new_n639_), .A2(new_n249_), .A3(new_n269_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n269_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT41), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n663_), .A3(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n647_), .B2(new_n432_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n432_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n639_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1327gat));
  NOR2_X1   g473(.A1(new_n587_), .A2(new_n646_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n457_), .A2(new_n458_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT103), .B1(new_n446_), .B2(new_n432_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n402_), .A2(new_n432_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n681_), .A2(new_n451_), .B1(new_n682_), .B2(new_n269_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n678_), .B1(new_n683_), .B2(new_n620_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n678_), .B(new_n620_), .C1(new_n449_), .C2(new_n461_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n675_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n675_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n450_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n643_), .A2(new_n646_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n588_), .A2(new_n693_), .ZN(new_n694_));
  OR3_X1    g493(.A1(new_n694_), .A2(G29gat), .A3(new_n450_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1328gat));
  NOR3_X1   g495(.A1(new_n694_), .A2(G36gat), .A3(new_n446_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT45), .Z(new_n698_));
  NAND4_X1  g497(.A1(new_n689_), .A2(KEYINPUT110), .A3(new_n655_), .A4(new_n690_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n655_), .A3(new_n690_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT111), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  AND4_X1   g503(.A1(KEYINPUT111), .A2(new_n703_), .A3(G36gat), .A4(new_n699_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT46), .B(new_n698_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  OAI21_X1  g509(.A(G43gat), .B1(new_n691_), .B2(new_n664_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n269_), .A2(new_n245_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n694_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT47), .Z(G1330gat));
  NAND4_X1  g513(.A1(new_n689_), .A2(G50gat), .A3(new_n672_), .A4(new_n690_), .ZN(new_n715_));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n694_), .B2(new_n432_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1331gat));
  NOR3_X1   g517(.A1(new_n462_), .A2(new_n548_), .A3(new_n586_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n637_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n375_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n548_), .A2(new_n636_), .A3(new_n586_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n645_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n450_), .A2(KEYINPUT112), .ZN(new_n726_));
  MUX2_X1   g525(.A(KEYINPUT112), .B(new_n726_), .S(G57gat), .Z(new_n727_));
  AOI21_X1  g526(.A(new_n722_), .B1(new_n725_), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n724_), .B2(new_n446_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n446_), .A2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n720_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n724_), .B2(new_n664_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n664_), .A2(G71gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n720_), .B2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n724_), .B2(new_n432_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n432_), .A2(G78gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n720_), .B2(new_n739_), .ZN(G1335gat));
  NAND2_X1  g539(.A1(new_n719_), .A2(new_n693_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n476_), .A3(new_n375_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n684_), .A2(new_n686_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n548_), .A2(new_n646_), .A3(new_n586_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT113), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n744_), .A2(new_n746_), .A3(new_n450_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(new_n476_), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n477_), .A3(new_n655_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n744_), .A2(new_n746_), .A3(new_n446_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n477_), .ZN(G1337gat));
  NOR2_X1   g550(.A1(new_n744_), .A2(new_n746_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n492_), .B1(new_n752_), .B2(new_n269_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n269_), .A2(new_n473_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n742_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g555(.A1(new_n742_), .A2(new_n474_), .A3(new_n672_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n752_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G106gat), .B1(new_n758_), .B2(new_n432_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g562(.A1(new_n586_), .A2(new_n636_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n619_), .A3(new_n548_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT118), .B1(new_n531_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n515_), .A2(new_n523_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n513_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT68), .B1(new_n775_), .B2(KEYINPUT12), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n527_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(KEYINPUT55), .A4(new_n525_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n525_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n778_), .A2(KEYINPUT117), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n773_), .A2(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n531_), .A2(new_n772_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n531_), .A2(KEYINPUT116), .A3(new_n772_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n785_), .A2(new_n790_), .A3(KEYINPUT119), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n542_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT119), .B1(new_n785_), .B2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n771_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n785_), .A2(new_n790_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n542_), .A4(new_n791_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n794_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n572_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n577_), .A2(new_n575_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n585_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n580_), .A2(new_n585_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n544_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n770_), .B1(new_n799_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n619_), .B1(new_n806_), .B2(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n586_), .A2(new_n544_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n803_), .A2(new_n802_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n643_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n643_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n808_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n769_), .B1(new_n817_), .B2(new_n636_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n375_), .B(new_n269_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT120), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n636_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT121), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(new_n825_), .A3(new_n636_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n769_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n586_), .B(new_n822_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G113gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n818_), .A2(new_n821_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n586_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n832_), .A2(G113gat), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(G1340gat));
  INV_X1    g634(.A(new_n548_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n822_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G120gat), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n831_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1341gat));
  OAI211_X1 g641(.A(new_n646_), .B(new_n822_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G127gat), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n832_), .A2(G127gat), .A3(new_n636_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1342gat));
  OAI211_X1 g645(.A(new_n620_), .B(new_n822_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G134gat), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n832_), .A2(G134gat), .A3(new_n643_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  NOR2_X1   g649(.A1(new_n269_), .A2(new_n432_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n823_), .B2(new_n768_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n655_), .A2(new_n450_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT122), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n856_));
  INV_X1    g655(.A(new_n854_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n818_), .A2(new_n856_), .A3(new_n852_), .A4(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n586_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G141gat), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n314_), .B(new_n586_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1344gat));
  OAI21_X1  g661(.A(new_n836_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G148gat), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n315_), .B(new_n836_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1345gat));
  OAI21_X1  g665(.A(new_n646_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n868_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n646_), .B(new_n870_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1346gat));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(new_n644_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n853_), .A2(new_n854_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n856_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n853_), .A2(KEYINPUT122), .A3(new_n854_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n619_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(new_n873_), .ZN(G1347gat));
  NAND3_X1  g678(.A1(new_n269_), .A2(new_n655_), .A3(new_n450_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n672_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n833_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G169gat), .B1(new_n827_), .B2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n827_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n883_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n886_), .ZN(new_n890_));
  OAI211_X1 g689(.A(G169gat), .B(new_n890_), .C1(new_n827_), .C2(new_n884_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(new_n889_), .A3(new_n891_), .ZN(G1348gat));
  NOR2_X1   g691(.A1(new_n827_), .A2(new_n882_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n836_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n818_), .A2(new_n672_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n548_), .A2(new_n214_), .A3(new_n880_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n214_), .B1(new_n895_), .B2(new_n896_), .ZN(G1349gat));
  NOR2_X1   g696(.A1(new_n880_), .A2(new_n636_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G183gat), .B1(new_n895_), .B2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n636_), .A2(new_n219_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n893_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n893_), .A2(new_n644_), .A3(new_n220_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n827_), .A2(new_n619_), .A3(new_n882_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n206_), .B2(new_n903_), .ZN(G1351gat));
  NOR2_X1   g703(.A1(new_n446_), .A2(new_n375_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n853_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n833_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT124), .B(G197gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1352gat));
  NAND3_X1  g708(.A1(new_n853_), .A2(new_n836_), .A3(new_n905_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n646_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n906_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT125), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n914_), .B(new_n916_), .ZN(G1354gat));
  NAND2_X1  g716(.A1(new_n620_), .A2(G218gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT127), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n906_), .A2(new_n919_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n853_), .A2(new_n644_), .A3(new_n905_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  AOI21_X1  g721(.A(G218gat), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n906_), .B2(new_n643_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n920_), .B1(new_n923_), .B2(new_n924_), .ZN(G1355gat));
endmodule


